magic
tech sky130A
magscale 1 2
timestamp 1687359403
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 842 2128 39546 597360
<< metal2 >>
rect 478 0 534 800
rect 846 0 902 800
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39486 0 39542 800
<< obsm2 >>
rect 478 856 39540 597349
rect 590 800 790 856
rect 958 800 1158 856
rect 1326 800 1526 856
rect 1694 800 1894 856
rect 2062 800 2262 856
rect 2430 800 2630 856
rect 2798 800 2998 856
rect 3166 800 3366 856
rect 3534 800 3734 856
rect 3902 800 4102 856
rect 4270 800 4470 856
rect 4638 800 4838 856
rect 5006 800 5206 856
rect 5374 800 5574 856
rect 5742 800 5942 856
rect 6110 800 6310 856
rect 6478 800 6678 856
rect 6846 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7782 856
rect 7950 800 8150 856
rect 8318 800 8518 856
rect 8686 800 8886 856
rect 9054 800 9254 856
rect 9422 800 9622 856
rect 9790 800 9990 856
rect 10158 800 10358 856
rect 10526 800 10726 856
rect 10894 800 11094 856
rect 11262 800 11462 856
rect 11630 800 11830 856
rect 11998 800 12198 856
rect 12366 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13302 856
rect 13470 800 13670 856
rect 13838 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16614 856
rect 16782 800 16982 856
rect 17150 800 17350 856
rect 17518 800 17718 856
rect 17886 800 18086 856
rect 18254 800 18454 856
rect 18622 800 18822 856
rect 18990 800 19190 856
rect 19358 800 19558 856
rect 19726 800 19926 856
rect 20094 800 20294 856
rect 20462 800 20662 856
rect 20830 800 21030 856
rect 21198 800 21398 856
rect 21566 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22502 856
rect 22670 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23606 856
rect 23774 800 23974 856
rect 24142 800 24342 856
rect 24510 800 24710 856
rect 24878 800 25078 856
rect 25246 800 25446 856
rect 25614 800 25814 856
rect 25982 800 26182 856
rect 26350 800 26550 856
rect 26718 800 26918 856
rect 27086 800 27286 856
rect 27454 800 27654 856
rect 27822 800 28022 856
rect 28190 800 28390 856
rect 28558 800 28758 856
rect 28926 800 29126 856
rect 29294 800 29494 856
rect 29662 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31334 856
rect 31502 800 31702 856
rect 31870 800 32070 856
rect 32238 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33174 856
rect 33342 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34646 856
rect 34814 800 35014 856
rect 35182 800 35382 856
rect 35550 800 35750 856
rect 35918 800 36118 856
rect 36286 800 36486 856
rect 36654 800 36854 856
rect 37022 800 37222 856
rect 37390 800 37590 856
rect 37758 800 37958 856
rect 38126 800 38326 856
rect 38494 800 38694 856
rect 38862 800 39062 856
rect 39230 800 39430 856
<< metal3 >>
rect 39200 584536 40000 584656
rect 0 573656 800 573776
rect 39200 559784 40000 559904
rect 39200 535032 40000 535152
rect 0 523880 800 524000
rect 39200 510280 40000 510400
rect 39200 485528 40000 485648
rect 0 474104 800 474224
rect 39200 460776 40000 460896
rect 39200 436024 40000 436144
rect 0 424328 800 424448
rect 39200 411272 40000 411392
rect 39200 386520 40000 386640
rect 0 374552 800 374672
rect 39200 361768 40000 361888
rect 39200 337016 40000 337136
rect 0 324776 800 324896
rect 39200 312264 40000 312384
rect 39200 287512 40000 287632
rect 0 275000 800 275120
rect 39200 262760 40000 262880
rect 39200 238008 40000 238128
rect 0 225224 800 225344
rect 39200 213256 40000 213376
rect 39200 188504 40000 188624
rect 0 175448 800 175568
rect 39200 163752 40000 163872
rect 39200 139000 40000 139120
rect 0 125672 800 125792
rect 39200 114248 40000 114368
rect 39200 89496 40000 89616
rect 0 75896 800 76016
rect 39200 64744 40000 64864
rect 39200 39992 40000 40112
rect 0 26120 800 26240
rect 39200 15240 40000 15360
<< obsm3 >>
rect 473 584736 39200 597345
rect 473 584456 39120 584736
rect 473 573856 39200 584456
rect 880 573576 39200 573856
rect 473 559984 39200 573576
rect 473 559704 39120 559984
rect 473 535232 39200 559704
rect 473 534952 39120 535232
rect 473 524080 39200 534952
rect 880 523800 39200 524080
rect 473 510480 39200 523800
rect 473 510200 39120 510480
rect 473 485728 39200 510200
rect 473 485448 39120 485728
rect 473 474304 39200 485448
rect 880 474024 39200 474304
rect 473 460976 39200 474024
rect 473 460696 39120 460976
rect 473 436224 39200 460696
rect 473 435944 39120 436224
rect 473 424528 39200 435944
rect 880 424248 39200 424528
rect 473 411472 39200 424248
rect 473 411192 39120 411472
rect 473 386720 39200 411192
rect 473 386440 39120 386720
rect 473 374752 39200 386440
rect 880 374472 39200 374752
rect 473 361968 39200 374472
rect 473 361688 39120 361968
rect 473 337216 39200 361688
rect 473 336936 39120 337216
rect 473 324976 39200 336936
rect 880 324696 39200 324976
rect 473 312464 39200 324696
rect 473 312184 39120 312464
rect 473 287712 39200 312184
rect 473 287432 39120 287712
rect 473 275200 39200 287432
rect 880 274920 39200 275200
rect 473 262960 39200 274920
rect 473 262680 39120 262960
rect 473 238208 39200 262680
rect 473 237928 39120 238208
rect 473 225424 39200 237928
rect 880 225144 39200 225424
rect 473 213456 39200 225144
rect 473 213176 39120 213456
rect 473 188704 39200 213176
rect 473 188424 39120 188704
rect 473 175648 39200 188424
rect 880 175368 39200 175648
rect 473 163952 39200 175368
rect 473 163672 39120 163952
rect 473 139200 39200 163672
rect 473 138920 39120 139200
rect 473 125872 39200 138920
rect 880 125592 39200 125872
rect 473 114448 39200 125592
rect 473 114168 39120 114448
rect 473 89696 39200 114168
rect 473 89416 39120 89696
rect 473 76096 39200 89416
rect 880 75816 39200 76096
rect 473 64944 39200 75816
rect 473 64664 39120 64944
rect 473 40192 39200 64664
rect 473 39912 39120 40192
rect 473 26320 39200 39912
rect 880 26040 39200 26320
rect 473 15440 39200 26040
rect 473 15160 39120 15440
rect 473 2143 39200 15160
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< obsm4 >>
rect 6683 2619 14477 24989
<< labels >>
rlabel metal3 s 39200 15240 40000 15360 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 275000 800 275120 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 89496 40000 89616 6 io_in[1]
port 4 nsew signal input
rlabel metal3 s 39200 163752 40000 163872 6 io_in[2]
port 5 nsew signal input
rlabel metal3 s 39200 238008 40000 238128 6 io_in[3]
port 6 nsew signal input
rlabel metal3 s 39200 312264 40000 312384 6 io_in[4]
port 7 nsew signal input
rlabel metal3 s 39200 386520 40000 386640 6 io_in[5]
port 8 nsew signal input
rlabel metal3 s 39200 460776 40000 460896 6 io_in[6]
port 9 nsew signal input
rlabel metal3 s 39200 535032 40000 535152 6 io_in[7]
port 10 nsew signal input
rlabel metal3 s 0 573656 800 573776 6 io_in[8]
port 11 nsew signal input
rlabel metal3 s 0 424328 800 424448 6 io_in[9]
port 12 nsew signal input
rlabel metal3 s 39200 64744 40000 64864 6 io_oeb[0]
port 13 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 io_oeb[10]
port 14 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[11]
port 15 nsew signal output
rlabel metal3 s 39200 139000 40000 139120 6 io_oeb[1]
port 16 nsew signal output
rlabel metal3 s 39200 213256 40000 213376 6 io_oeb[2]
port 17 nsew signal output
rlabel metal3 s 39200 287512 40000 287632 6 io_oeb[3]
port 18 nsew signal output
rlabel metal3 s 39200 361768 40000 361888 6 io_oeb[4]
port 19 nsew signal output
rlabel metal3 s 39200 436024 40000 436144 6 io_oeb[5]
port 20 nsew signal output
rlabel metal3 s 39200 510280 40000 510400 6 io_oeb[6]
port 21 nsew signal output
rlabel metal3 s 39200 584536 40000 584656 6 io_oeb[7]
port 22 nsew signal output
rlabel metal3 s 0 474104 800 474224 6 io_oeb[8]
port 23 nsew signal output
rlabel metal3 s 0 324776 800 324896 6 io_oeb[9]
port 24 nsew signal output
rlabel metal3 s 39200 39992 40000 40112 6 io_out[0]
port 25 nsew signal output
rlabel metal3 s 0 225224 800 225344 6 io_out[10]
port 26 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 io_out[11]
port 27 nsew signal output
rlabel metal3 s 39200 114248 40000 114368 6 io_out[1]
port 28 nsew signal output
rlabel metal3 s 39200 188504 40000 188624 6 io_out[2]
port 29 nsew signal output
rlabel metal3 s 39200 262760 40000 262880 6 io_out[3]
port 30 nsew signal output
rlabel metal3 s 39200 337016 40000 337136 6 io_out[4]
port 31 nsew signal output
rlabel metal3 s 39200 411272 40000 411392 6 io_out[5]
port 32 nsew signal output
rlabel metal3 s 39200 485528 40000 485648 6 io_out[6]
port 33 nsew signal output
rlabel metal3 s 39200 559784 40000 559904 6 io_out[7]
port 34 nsew signal output
rlabel metal3 s 0 523880 800 524000 6 io_out[8]
port 35 nsew signal output
rlabel metal3 s 0 374552 800 374672 6 io_out[9]
port 36 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 irq
port 37 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 38 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 38 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 39 nsew ground bidirectional
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 40 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 41 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 42 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_adr_i[0]
port 43 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[10]
port 44 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[11]
port 45 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[12]
port 46 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[13]
port 47 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[14]
port 48 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[15]
port 49 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[16]
port 50 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[17]
port 51 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_adr_i[18]
port 52 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[19]
port 53 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[1]
port 54 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[20]
port 55 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[21]
port 56 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_adr_i[22]
port 57 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[23]
port 58 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[24]
port 59 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_adr_i[25]
port 60 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[26]
port 61 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[27]
port 62 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_adr_i[28]
port 63 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[29]
port 64 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[2]
port 65 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[30]
port 66 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_adr_i[31]
port 67 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[3]
port 68 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[4]
port 69 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[5]
port 70 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[6]
port 71 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[7]
port 72 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[8]
port 73 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[9]
port 74 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_cyc_i
port 75 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[0]
port 76 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[10]
port 77 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[11]
port 78 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[12]
port 79 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[13]
port 80 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[14]
port 81 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[15]
port 82 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[16]
port 83 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[17]
port 84 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[18]
port 85 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[19]
port 86 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[1]
port 87 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[20]
port 88 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[21]
port 89 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[22]
port 90 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[23]
port 91 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[24]
port 92 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[25]
port 93 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[26]
port 94 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[27]
port 95 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_i[28]
port 96 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[29]
port 97 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[2]
port 98 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[30]
port 99 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[31]
port 100 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[3]
port 101 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[4]
port 102 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[5]
port 103 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[6]
port 104 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[7]
port 105 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[8]
port 106 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[9]
port 107 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 108 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[10]
port 109 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[11]
port 110 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[12]
port 111 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[13]
port 112 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[14]
port 113 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[15]
port 114 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[16]
port 115 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[17]
port 116 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_o[18]
port 117 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[19]
port 118 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[1]
port 119 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[20]
port 120 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[21]
port 121 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[22]
port 122 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[23]
port 123 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[24]
port 124 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[25]
port 125 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[26]
port 126 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[27]
port 127 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[28]
port 128 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[29]
port 129 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[2]
port 130 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[30]
port 131 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[31]
port 132 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[3]
port 133 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_o[4]
port 134 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[5]
port 135 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[6]
port 136 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[7]
port 137 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[8]
port 138 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[9]
port 139 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 140 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_sel_i[1]
port 141 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_sel_i[2]
port 142 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_sel_i[3]
port 143 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_stb_i
port 144 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_we_i
port 145 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8209004
string GDS_FILE /home/hosni/OpenLane-tutorial/7-segment/openlane/user_proj_example2/runs/23_06_21_07_54/results/signoff/user_proj_example2.magic.gds
string GDS_START 591128
<< end >>


// This is the unpowered netlist.
module user_proj_example1 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [11:0] io_in;
 output [11:0] io_oeb;
 output [11:0] io_out;

 wire net25;
 wire net35;
 wire net36;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net37;
 wire \Clock_part1.dig_cnt[0] ;
 wire \Clock_part1.dig_cnt[1] ;
 wire \Clock_part1.min_ones[0] ;
 wire \Clock_part1.min_ones[1] ;
 wire \Clock_part1.min_ones[2] ;
 wire \Clock_part1.min_ones[3] ;
 wire \Clock_part1.min_tens[0] ;
 wire \Clock_part1.min_tens[1] ;
 wire \Clock_part1.min_tens[2] ;
 wire \Clock_part1.min_tens[3] ;
 wire \Clock_part1.scan ;
 wire \Clock_part1.scan_div[0] ;
 wire \Clock_part1.scan_div[10] ;
 wire \Clock_part1.scan_div[11] ;
 wire \Clock_part1.scan_div[12] ;
 wire \Clock_part1.scan_div[13] ;
 wire \Clock_part1.scan_div[14] ;
 wire \Clock_part1.scan_div[15] ;
 wire \Clock_part1.scan_div[16] ;
 wire \Clock_part1.scan_div[17] ;
 wire \Clock_part1.scan_div[18] ;
 wire \Clock_part1.scan_div[19] ;
 wire \Clock_part1.scan_div[1] ;
 wire \Clock_part1.scan_div[20] ;
 wire \Clock_part1.scan_div[21] ;
 wire \Clock_part1.scan_div[22] ;
 wire \Clock_part1.scan_div[23] ;
 wire \Clock_part1.scan_div[24] ;
 wire \Clock_part1.scan_div[25] ;
 wire \Clock_part1.scan_div[26] ;
 wire \Clock_part1.scan_div[27] ;
 wire \Clock_part1.scan_div[28] ;
 wire \Clock_part1.scan_div[29] ;
 wire \Clock_part1.scan_div[2] ;
 wire \Clock_part1.scan_div[30] ;
 wire \Clock_part1.scan_div[31] ;
 wire \Clock_part1.scan_div[3] ;
 wire \Clock_part1.scan_div[4] ;
 wire \Clock_part1.scan_div[5] ;
 wire \Clock_part1.scan_div[6] ;
 wire \Clock_part1.scan_div[7] ;
 wire \Clock_part1.scan_div[8] ;
 wire \Clock_part1.scan_div[9] ;
 wire \Clock_part1.sec ;
 wire \Clock_part1.sec_div[0] ;
 wire \Clock_part1.sec_div[10] ;
 wire \Clock_part1.sec_div[11] ;
 wire \Clock_part1.sec_div[12] ;
 wire \Clock_part1.sec_div[13] ;
 wire \Clock_part1.sec_div[14] ;
 wire \Clock_part1.sec_div[15] ;
 wire \Clock_part1.sec_div[16] ;
 wire \Clock_part1.sec_div[17] ;
 wire \Clock_part1.sec_div[18] ;
 wire \Clock_part1.sec_div[19] ;
 wire \Clock_part1.sec_div[1] ;
 wire \Clock_part1.sec_div[20] ;
 wire \Clock_part1.sec_div[21] ;
 wire \Clock_part1.sec_div[22] ;
 wire \Clock_part1.sec_div[23] ;
 wire \Clock_part1.sec_div[24] ;
 wire \Clock_part1.sec_div[25] ;
 wire \Clock_part1.sec_div[26] ;
 wire \Clock_part1.sec_div[27] ;
 wire \Clock_part1.sec_div[28] ;
 wire \Clock_part1.sec_div[29] ;
 wire \Clock_part1.sec_div[2] ;
 wire \Clock_part1.sec_div[30] ;
 wire \Clock_part1.sec_div[31] ;
 wire \Clock_part1.sec_div[3] ;
 wire \Clock_part1.sec_div[4] ;
 wire \Clock_part1.sec_div[5] ;
 wire \Clock_part1.sec_div[6] ;
 wire \Clock_part1.sec_div[7] ;
 wire \Clock_part1.sec_div[8] ;
 wire \Clock_part1.sec_div[9] ;
 wire \Clock_part1.sec_ones[0] ;
 wire \Clock_part1.sec_ones[1] ;
 wire \Clock_part1.sec_ones[2] ;
 wire \Clock_part1.sec_ones[3] ;
 wire \Clock_part1.sec_tens[0] ;
 wire \Clock_part1.sec_tens[1] ;
 wire \Clock_part1.sec_tens[2] ;
 wire \Clock_part1.sec_tens[3] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_213_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_209_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_209_));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1000_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1000_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1000_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1001_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1001_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1001_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1001_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1001_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1002_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1002_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1002_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1003_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1003_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1003_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1003_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1003_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1004_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1004_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1004_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1005_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1005_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1005_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1005_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1005_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1006_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1006_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1006_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1007_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1007_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1007_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1007_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1007_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1008_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1008_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1008_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1009_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1009_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1009_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1009_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1009_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1010_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1010_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1010_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1011_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1011_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1011_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1011_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1011_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1012_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1012_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1012_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1013_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1013_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1013_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1013_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1013_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1014_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1014_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1014_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1015_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1015_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1015_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1015_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1015_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1016_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1016_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1016_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1017_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1017_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1017_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1017_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1017_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1018_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1018_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1018_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1019_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1019_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1019_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1019_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1019_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1020_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1020_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1020_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1021_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1021_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1021_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1021_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1021_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1022_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1022_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1022_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1023_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1023_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1023_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1023_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1023_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1024_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1024_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1024_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1025_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1025_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1025_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1025_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1025_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1026_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1026_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1026_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1027_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1027_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1027_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1027_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1027_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_1028_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1028_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1028_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1028_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1029_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1029_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1029_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1029_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1029_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1030_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1030_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1030_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1031_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1031_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1031_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1031_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1031_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1032_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1032_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1032_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1033_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1033_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1033_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1033_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1033_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1034_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1034_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1034_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1035_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1035_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1035_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1035_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1035_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1036_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1036_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1036_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1037_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1037_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1037_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1037_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1037_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1038_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1038_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1038_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1039_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1039_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1039_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1039_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1039_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1040_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1040_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1040_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1041_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1041_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1041_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1041_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1041_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1042_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1042_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1042_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1043_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1043_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1043_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1043_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1043_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1044_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1044_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1044_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1045_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1045_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1045_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1045_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1045_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1046_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1046_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1046_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1047_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1047_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1047_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1047_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1047_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1048_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1048_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1048_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1049_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1049_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1049_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1049_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1049_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1050_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1050_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1050_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1051_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1051_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1051_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1051_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1051_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1052_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1052_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1052_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1053_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1053_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1053_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1053_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1053_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1054_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1054_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1054_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1055_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1055_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1055_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1055_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1055_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1056_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1056_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1056_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1057_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1057_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1057_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1057_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1057_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1058_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1058_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1058_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1059_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1059_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1059_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1059_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1059_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1060_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1060_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1060_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1061_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1061_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1061_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1061_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1061_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1062_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1062_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1062_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1063_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1063_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1063_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1063_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1063_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1064_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1064_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1064_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1065_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1065_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1065_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1065_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1065_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1066_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1066_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1066_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1067_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1067_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1067_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1067_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1067_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1068_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1068_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1068_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1069_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1069_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1069_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1069_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1069_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1070_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1070_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1070_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1071_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1071_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1071_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1071_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1071_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1072_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1072_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1072_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1073_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1073_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1073_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1073_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1073_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_1074_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1074_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1074_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1074_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1075_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1075_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1075_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1075_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1075_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1076_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1076_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1076_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1077_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1077_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1077_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1077_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1077_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1078_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1078_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1078_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1079_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1079_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1079_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1079_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1079_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1080_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1080_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1080_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1081_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1081_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1081_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1081_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1081_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1082_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1082_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1082_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1083_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1083_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1083_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1083_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1083_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1084_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1084_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1084_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1085_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1085_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1085_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1085_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1085_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1086_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1086_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1086_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1087_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1087_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1087_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1087_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1087_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1088_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1088_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1088_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1089_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1089_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1089_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1089_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1089_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1090_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1090_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1090_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1091_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1091_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1091_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1091_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1091_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1092_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1092_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1092_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1093_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1093_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_1093_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1093_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_286_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_287_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_287_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_287_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_288_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_289_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_289_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_289_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_290_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_291_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_291_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_291_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_293_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_293_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_293_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_293_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_294_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_295_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_295_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_295_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_296_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_297_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_297_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_297_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_297_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_298_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_299_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_299_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_300_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_301_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_301_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_301_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_301_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_302_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_303_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_303_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_303_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_303_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_304_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_305_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_305_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_305_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_305_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_306_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_307_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_307_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_307_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_307_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_307_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_308_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_309_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_309_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_309_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_309_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_311_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_311_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_311_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_311_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_312_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_313_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_313_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_313_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_313_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_314_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_315_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_315_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_315_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_315_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_317_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_317_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_317_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_317_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_318_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_318_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_318_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_318_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_319_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_319_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_319_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_320_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_321_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_321_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_321_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_321_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_321_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_322_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_322_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_322_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_323_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_323_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_323_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_323_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_323_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_324_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_324_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_325_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_325_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_325_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_325_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_326_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_327_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_327_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_327_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_327_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_328_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_329_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_329_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_329_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_329_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_329_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_330_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_331_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_331_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_331_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_331_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_331_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_332_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_333_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_333_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_333_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_333_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_333_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_335_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_335_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_335_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_335_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_335_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_337_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_337_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_337_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_337_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_337_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_338_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_339_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_339_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_339_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_339_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_339_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_340_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_340_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_340_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_341_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_341_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_341_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_341_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_342_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_342_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_342_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_342_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_343_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_343_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_343_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_343_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_343_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_344_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_345_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_345_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_345_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_345_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_345_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_346_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_347_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_347_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_347_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_347_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_347_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_348_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_349_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_349_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_349_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_349_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_349_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_350_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_351_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_351_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_351_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_351_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_351_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_352_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_353_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_353_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_353_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_353_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_353_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_355_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_355_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_355_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_355_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_356_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_357_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_357_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_357_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_357_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_358_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_358_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_358_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_359_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_359_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_359_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_359_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_359_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_360_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_360_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_360_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_361_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_361_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_361_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_361_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_361_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_362_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_362_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_362_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_363_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_363_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_363_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_363_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_363_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_364_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_364_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_364_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_365_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_365_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_365_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_365_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_365_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_366_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_366_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_366_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_367_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_367_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_367_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_367_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_367_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_368_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_368_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_368_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_369_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_369_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_369_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_369_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_369_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_370_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_370_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_370_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_371_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_371_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_371_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_371_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_371_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_372_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_372_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_372_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_373_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_373_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_373_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_373_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_373_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_374_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_374_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_374_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_375_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_375_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_375_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_375_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_375_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_376_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_376_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_376_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_377_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_377_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_377_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_377_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_377_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_378_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_378_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_378_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_379_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_379_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_379_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_379_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_379_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_380_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_380_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_380_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_381_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_381_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_381_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_381_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_381_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_382_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_382_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_382_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_383_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_383_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_383_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_383_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_383_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_384_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_384_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_384_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_385_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_385_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_385_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_385_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_385_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_386_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_386_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_386_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_387_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_387_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_387_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_387_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_387_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_387_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_388_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_388_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_388_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_389_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_389_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_389_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_389_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_389_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_390_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_390_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_390_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_391_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_391_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_391_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_391_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_391_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_392_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_392_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_392_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_393_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_393_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_393_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_393_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_393_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_394_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_394_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_394_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_395_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_395_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_395_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_395_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_395_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_396_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_396_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_396_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_397_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_397_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_397_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_397_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_397_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_398_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_398_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_398_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_399_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_399_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_399_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_399_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_399_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_400_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_400_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_400_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_401_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_401_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_401_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_401_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_401_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_402_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_402_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_402_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_403_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_403_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_403_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_403_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_403_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_404_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_404_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_404_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_405_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_405_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_405_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_405_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_405_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_406_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_406_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_406_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_407_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_407_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_407_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_407_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_407_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_408_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_408_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_408_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_409_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_409_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_409_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_409_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_409_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_410_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_410_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_410_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_410_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_411_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_411_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_411_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_411_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_411_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_412_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_412_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_412_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_413_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_413_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_413_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_413_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_413_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_414_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_414_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_414_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_415_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_415_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_415_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_415_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_415_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_416_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_416_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_416_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_417_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_417_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_417_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_417_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_417_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_418_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_418_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_418_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_419_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_419_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_419_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_419_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_419_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_420_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_420_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_420_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_421_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_421_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_421_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_421_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_421_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_422_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_422_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_422_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_423_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_423_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_423_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_423_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_423_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_424_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_424_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_424_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_425_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_425_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_425_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_425_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_425_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_426_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_426_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_426_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_427_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_427_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_427_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_427_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_427_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_428_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_428_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_428_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_429_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_429_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_429_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_429_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_429_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_430_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_430_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_430_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_431_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_431_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_431_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_431_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_431_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_432_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_432_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_432_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_433_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_433_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_433_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_433_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_433_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_434_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_434_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_434_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_435_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_435_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_435_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_435_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_435_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_436_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_436_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_436_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_437_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_437_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_437_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_437_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_437_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_438_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_438_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_438_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_439_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_439_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_439_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_439_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_439_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_440_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_440_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_440_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_441_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_441_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_441_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_441_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_441_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_442_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_442_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_442_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_443_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_443_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_443_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_443_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_443_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_444_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_444_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_444_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_445_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_445_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_445_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_445_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_445_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_446_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_446_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_446_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_447_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_447_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_447_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_447_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_447_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_448_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_448_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_448_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_449_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_449_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_449_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_449_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_449_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_450_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_450_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_450_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_451_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_451_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_451_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_451_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_451_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_452_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_452_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_452_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_453_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_453_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_453_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_453_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_453_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_454_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_454_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_454_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_455_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_455_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_455_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_455_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_455_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_456_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_456_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_456_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_457_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_457_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_457_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_457_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_457_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_458_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_458_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_458_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_459_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_459_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_459_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_459_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_459_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_460_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_460_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_460_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_461_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_461_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_461_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_461_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_461_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_462_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_462_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_462_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_463_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_463_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_463_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_463_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_463_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_464_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_464_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_464_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_465_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_465_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_465_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_465_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_465_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_466_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_466_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_466_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_467_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_467_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_467_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_467_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_467_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_468_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_468_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_468_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_469_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_469_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_469_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_469_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_469_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_470_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_470_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_470_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_471_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_471_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_471_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_471_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_471_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_472_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_472_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_472_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_473_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_473_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_473_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_473_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_473_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_474_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_474_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_474_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_475_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_475_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_475_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_475_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_475_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_476_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_476_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_476_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_477_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_477_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_477_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_477_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_477_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_478_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_478_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_478_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_478_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_478_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_478_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_479_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_479_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_479_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_479_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_479_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_480_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_480_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_480_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_481_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_481_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_481_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_481_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_481_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_482_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_482_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_482_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_483_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_483_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_483_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_483_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_483_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_484_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_484_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_484_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_485_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_485_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_485_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_485_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_485_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_486_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_486_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_486_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_487_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_487_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_487_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_487_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_487_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_488_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_488_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_488_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_489_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_489_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_489_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_489_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_489_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_490_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_490_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_490_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_491_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_491_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_491_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_491_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_491_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_492_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_492_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_492_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_493_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_493_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_493_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_493_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_493_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_494_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_494_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_494_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_495_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_495_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_495_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_495_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_495_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_496_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_496_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_496_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_497_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_497_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_497_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_497_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_497_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_498_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_498_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_498_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_499_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_499_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_499_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_499_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_499_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_500_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_500_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_500_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_501_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_501_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_501_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_501_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_501_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_502_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_502_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_502_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_503_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_503_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_503_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_503_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_503_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_504_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_504_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_504_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_505_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_505_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_505_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_505_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_505_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_506_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_506_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_506_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_507_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_507_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_507_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_507_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_507_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_508_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_508_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_508_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_509_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_509_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_509_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_509_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_509_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_510_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_510_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_510_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_511_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_511_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_511_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_511_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_511_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_512_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_512_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_512_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_513_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_513_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_513_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_513_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_513_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_514_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_514_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_514_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_515_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_515_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_515_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_515_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_515_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_516_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_516_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_516_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_517_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_517_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_517_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_517_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_517_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_518_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_518_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_518_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_519_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_519_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_519_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_519_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_519_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_520_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_520_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_520_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_521_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_521_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_521_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_521_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_521_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_522_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_522_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_522_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_523_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_523_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_523_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_523_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_523_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_524_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_524_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_524_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_525_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_525_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_525_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_525_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_525_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_525_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_526_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_526_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_526_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_527_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_527_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_527_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_527_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_527_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_528_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_528_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_528_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_529_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_529_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_529_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_529_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_529_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_530_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_530_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_530_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_531_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_531_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_531_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_531_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_531_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_532_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_532_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_532_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_533_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_533_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_533_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_533_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_533_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_534_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_534_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_534_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_535_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_535_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_535_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_535_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_535_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_536_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_536_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_536_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_537_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_537_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_537_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_537_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_537_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_538_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_538_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_538_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_539_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_539_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_539_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_539_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_539_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_540_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_540_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_540_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_541_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_541_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_541_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_541_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_541_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_542_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_542_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_542_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_543_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_543_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_543_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_543_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_543_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_544_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_544_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_544_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_545_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_545_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_545_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_545_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_545_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_546_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_546_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_546_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_547_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_547_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_547_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_547_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_547_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_548_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_548_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_548_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_549_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_549_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_549_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_549_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_549_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_550_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_550_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_550_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_551_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_551_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_551_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_551_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_551_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_552_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_552_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_552_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_553_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_553_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_553_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_553_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_553_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_554_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_554_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_554_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_555_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_555_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_555_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_555_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_555_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_556_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_556_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_556_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_557_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_557_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_557_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_557_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_557_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_558_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_558_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_558_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_559_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_559_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_559_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_559_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_559_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_560_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_560_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_560_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_561_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_561_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_561_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_561_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_561_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_562_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_562_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_562_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_563_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_563_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_563_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_563_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_563_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_564_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_564_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_564_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_565_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_565_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_565_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_565_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_565_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_566_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_566_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_566_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_567_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_567_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_567_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_567_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_567_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_568_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_568_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_568_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_569_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_569_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_569_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_569_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_569_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_570_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_570_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_570_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_571_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_571_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_571_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_571_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_571_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_572_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_572_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_572_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_573_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_573_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_573_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_573_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_573_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_574_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_574_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_574_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_575_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_575_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_575_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_575_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_575_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_576_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_576_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_576_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_577_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_577_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_577_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_577_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_577_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_578_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_578_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_578_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_579_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_579_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_579_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_579_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_579_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_580_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_580_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_580_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_581_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_581_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_581_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_581_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_581_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_582_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_582_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_582_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_583_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_583_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_583_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_583_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_583_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_584_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_584_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_584_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_585_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_585_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_585_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_585_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_585_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_586_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_586_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_586_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_587_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_587_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_587_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_587_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_587_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_588_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_588_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_588_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_589_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_589_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_589_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_589_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_589_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_590_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_590_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_590_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_591_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_591_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_591_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_591_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_591_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_592_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_592_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_592_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_593_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_593_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_593_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_593_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_594_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_594_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_594_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_595_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_595_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_595_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_595_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_595_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_596_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_596_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_596_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_597_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_597_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_597_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_597_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_597_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_598_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_598_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_598_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_599_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_599_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_599_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_599_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_599_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_600_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_600_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_600_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_601_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_601_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_601_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_601_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_601_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_602_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_602_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_602_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_603_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_603_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_603_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_603_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_603_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_604_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_604_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_604_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_605_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_605_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_605_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_605_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_605_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_606_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_606_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_606_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_607_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_607_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_607_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_607_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_607_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_608_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_608_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_608_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_609_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_609_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_609_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_609_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_609_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_610_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_610_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_610_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_611_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_611_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_611_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_611_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_611_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_612_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_612_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_612_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_613_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_613_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_613_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_613_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_613_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_613_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_614_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_614_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_614_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_614_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_614_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_615_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_615_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_615_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_615_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_615_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_615_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_615_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_615_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_616_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_616_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_616_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_616_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_616_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_617_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_617_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_617_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_617_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_617_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_617_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_617_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_617_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_618_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_618_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_618_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_618_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_618_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_618_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_619_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_619_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_619_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_619_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_619_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_619_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_620_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_620_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_620_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_621_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_621_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_621_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_621_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_621_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_622_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_622_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_622_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_623_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_623_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_623_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_623_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_623_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_624_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_624_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_624_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_625_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_625_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_625_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_625_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_625_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_626_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_626_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_626_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_627_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_627_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_627_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_627_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_627_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_628_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_628_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_628_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_629_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_629_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_629_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_629_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_629_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_630_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_630_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_630_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_631_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_631_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_631_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_631_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_631_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_632_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_632_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_632_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_633_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_633_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_633_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_633_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_633_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_634_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_634_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_634_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_635_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_635_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_635_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_635_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_635_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_636_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_636_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_636_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_637_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_637_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_637_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_637_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_637_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_638_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_638_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_638_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_639_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_639_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_639_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_639_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_639_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_640_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_640_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_640_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_641_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_641_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_641_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_641_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_641_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_642_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_642_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_642_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_643_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_643_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_643_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_643_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_643_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_644_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_644_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_644_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_645_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_645_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_645_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_645_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_645_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_646_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_646_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_646_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_647_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_647_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_647_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_647_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_647_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_648_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_648_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_648_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_649_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_649_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_649_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_649_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_649_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_650_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_650_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_650_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_651_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_651_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_651_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_651_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_651_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_652_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_652_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_652_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_653_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_653_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_653_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_653_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_653_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_654_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_654_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_654_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_655_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_655_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_655_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_655_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_655_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_656_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_656_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_656_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_657_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_657_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_657_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_657_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_657_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_658_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_658_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_658_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_659_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_659_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_659_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_659_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_659_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_660_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_660_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_660_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_661_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_661_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_661_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_661_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_661_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_662_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_662_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_662_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_662_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_663_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_663_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_663_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_663_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_663_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_664_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_664_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_664_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_665_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_665_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_665_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_665_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_665_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_666_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_666_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_666_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_667_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_667_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_667_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_667_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_667_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_668_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_668_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_668_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_669_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_669_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_669_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_669_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_669_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_670_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_670_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_670_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_671_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_671_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_671_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_671_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_671_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_672_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_672_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_672_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_673_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_673_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_673_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_673_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_673_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_674_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_674_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_674_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_675_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_675_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_675_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_675_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_675_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_676_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_676_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_676_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_677_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_677_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_677_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_677_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_677_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_678_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_678_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_678_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_679_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_679_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_679_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_679_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_679_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_680_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_680_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_680_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_681_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_681_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_681_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_681_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_681_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_682_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_682_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_682_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_683_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_683_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_683_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_683_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_683_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_684_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_684_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_684_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_685_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_685_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_685_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_685_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_685_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_685_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_685_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_686_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_686_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_686_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_687_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_687_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_687_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_687_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_687_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_688_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_688_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_688_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_689_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_689_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_689_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_689_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_689_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_690_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_690_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_690_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_691_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_691_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_691_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_691_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_691_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_692_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_692_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_692_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_693_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_693_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_693_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_693_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_693_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_694_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_694_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_694_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_695_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_695_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_695_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_695_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_695_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_696_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_696_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_696_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_697_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_697_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_697_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_697_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_697_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_698_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_698_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_698_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_699_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_699_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_699_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_699_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_699_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_700_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_700_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_700_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_701_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_701_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_701_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_701_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_701_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_702_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_702_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_702_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_703_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_703_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_703_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_703_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_703_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_704_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_704_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_704_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_705_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_705_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_705_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_705_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_705_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_706_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_706_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_706_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_707_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_707_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_707_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_707_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_707_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_708_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_708_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_708_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_709_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_709_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_709_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_709_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_709_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_710_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_710_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_710_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_711_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_711_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_711_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_711_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_711_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_712_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_712_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_712_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_713_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_713_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_713_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_713_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_713_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_714_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_714_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_714_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_715_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_715_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_715_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_715_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_715_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_716_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_716_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_716_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_717_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_717_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_717_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_717_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_717_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_718_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_718_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_718_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_719_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_719_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_719_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_719_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_719_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_720_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_720_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_720_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_721_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_721_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_721_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_721_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_721_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_722_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_722_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_722_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_723_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_723_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_723_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_723_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_723_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_724_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_724_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_724_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_725_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_725_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_725_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_725_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_725_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_726_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_726_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_726_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_727_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_727_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_727_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_727_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_727_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_728_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_728_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_728_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_729_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_729_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_729_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_729_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_729_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_730_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_730_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_730_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_731_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_731_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_731_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_731_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_731_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_732_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_732_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_732_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_733_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_733_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_733_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_733_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_733_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_734_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_734_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_734_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_735_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_735_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_735_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_735_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_735_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_736_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_736_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_736_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_737_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_737_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_737_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_737_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_737_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_738_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_738_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_738_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_739_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_739_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_739_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_739_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_739_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_740_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_740_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_740_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_741_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_741_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_741_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_741_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_741_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_742_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_742_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_742_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_743_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_743_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_743_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_743_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_743_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_744_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_744_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_744_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_745_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_745_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_745_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_745_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_745_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_746_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_746_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_746_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_747_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_747_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_747_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_747_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_747_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_748_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_748_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_748_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_749_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_749_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_749_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_749_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_749_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_750_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_750_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_750_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_751_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_751_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_751_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_751_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_751_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_752_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_752_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_752_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_752_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_753_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_753_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_753_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_753_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_753_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_754_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_754_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_754_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_755_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_755_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_755_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_755_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_755_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_756_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_756_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_756_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_757_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_757_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_757_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_757_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_757_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_758_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_758_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_758_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_759_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_759_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_759_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_759_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_759_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_760_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_760_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_760_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_761_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_761_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_761_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_761_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_761_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_762_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_762_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_762_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_763_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_763_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_763_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_763_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_763_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_764_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_764_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_764_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_765_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_765_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_765_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_765_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_765_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_766_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_766_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_766_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_767_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_767_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_767_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_767_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_767_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_768_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_768_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_768_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_769_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_769_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_769_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_769_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_769_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_770_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_770_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_770_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_771_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_771_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_771_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_771_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_771_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_772_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_772_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_772_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_773_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_773_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_773_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_773_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_773_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_774_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_774_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_774_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_775_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_775_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_775_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_775_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_775_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_776_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_776_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_776_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_777_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_777_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_777_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_777_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_777_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_778_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_778_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_778_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_779_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_779_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_779_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_779_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_779_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_780_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_780_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_780_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_781_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_781_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_781_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_781_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_781_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_782_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_782_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_782_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_783_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_783_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_783_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_783_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_783_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_784_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_784_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_784_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_785_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_785_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_785_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_785_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_785_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_786_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_786_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_786_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_787_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_787_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_787_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_787_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_787_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_788_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_788_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_788_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_789_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_789_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_789_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_789_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_789_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_790_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_790_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_790_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_791_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_791_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_791_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_791_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_791_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_792_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_792_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_792_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_793_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_793_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_793_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_793_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_793_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_794_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_794_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_794_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_795_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_795_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_795_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_795_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_795_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_796_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_796_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_796_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_797_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_797_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_797_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_797_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_797_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_798_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_798_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_798_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_799_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_799_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_799_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_799_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_799_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_799_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_800_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_800_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_800_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_801_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_801_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_801_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_801_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_801_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_802_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_802_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_802_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_803_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_803_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_803_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_803_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_803_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_804_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_804_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_804_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_805_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_805_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_805_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_805_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_805_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_806_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_806_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_806_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_807_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_807_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_807_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_807_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_807_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_808_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_808_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_808_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_809_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_809_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_809_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_809_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_809_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_810_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_810_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_810_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_811_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_811_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_811_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_811_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_811_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_812_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_812_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_812_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_813_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_813_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_813_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_813_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_813_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_814_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_814_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_814_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_815_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_815_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_815_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_815_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_815_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_816_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_816_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_816_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_817_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_817_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_817_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_817_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_817_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_818_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_818_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_818_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_819_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_819_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_819_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_819_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_819_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_820_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_820_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_820_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_821_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_821_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_821_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_821_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_821_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_822_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_822_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_822_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_823_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_823_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_823_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_823_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_823_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_824_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_824_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_824_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_825_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_825_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_825_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_825_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_825_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_826_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_826_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_826_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_827_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_827_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_827_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_827_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_827_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_828_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_828_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_828_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_829_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_829_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_829_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_829_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_829_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_830_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_830_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_830_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_831_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_831_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_831_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_831_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_831_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_832_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_832_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_832_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_833_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_833_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_833_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_833_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_833_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_834_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_834_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_834_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_835_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_835_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_835_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_835_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_835_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_836_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_836_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_836_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_837_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_837_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_837_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_837_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_837_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_838_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_838_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_838_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_839_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_839_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_839_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_839_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_839_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_840_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_840_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_840_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_841_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_841_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_841_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_841_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_841_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_842_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_842_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_842_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_843_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_843_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_843_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_843_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_843_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_844_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_844_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_844_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_845_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_845_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_845_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_845_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_845_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_846_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_846_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_846_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_847_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_847_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_847_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_847_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_847_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_848_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_848_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_848_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_849_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_849_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_849_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_849_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_849_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_850_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_850_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_850_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_851_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_851_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_851_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_851_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_851_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_852_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_852_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_852_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_853_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_853_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_853_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_853_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_853_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_854_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_854_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_854_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_855_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_855_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_855_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_855_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_855_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_856_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_856_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_856_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_857_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_857_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_857_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_857_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_857_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_858_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_858_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_858_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_859_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_859_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_859_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_859_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_859_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_860_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_860_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_860_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_861_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_861_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_861_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_861_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_861_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_862_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_862_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_862_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_863_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_863_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_863_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_863_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_863_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_864_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_864_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_864_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_865_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_865_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_865_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_865_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_865_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_866_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_866_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_866_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_867_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_867_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_867_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_867_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_867_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_868_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_868_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_868_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_869_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_869_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_869_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_869_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_869_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_870_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_870_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_870_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_871_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_871_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_871_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_871_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_871_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_872_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_872_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_872_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_873_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_873_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_873_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_873_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_873_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_874_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_874_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_874_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_875_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_875_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_875_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_875_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_875_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_876_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_876_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_876_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_877_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_877_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_877_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_877_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_877_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_878_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_878_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_878_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_879_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_879_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_879_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_879_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_879_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_880_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_880_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_880_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_881_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_881_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_881_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_881_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_881_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_882_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_882_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_882_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_883_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_883_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_883_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_883_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_883_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_884_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_884_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_884_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_885_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_885_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_885_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_885_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_885_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_886_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_886_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_886_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_887_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_887_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_887_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_887_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_887_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_888_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_888_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_888_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_889_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_889_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_889_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_889_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_889_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_890_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_890_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_890_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_890_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_891_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_891_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_891_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_891_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_891_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_892_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_892_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_892_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_893_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_893_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_893_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_893_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_893_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_894_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_894_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_894_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_895_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_895_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_895_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_895_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_895_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_896_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_896_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_896_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_897_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_897_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_897_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_897_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_897_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_898_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_898_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_898_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_899_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_899_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_899_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_899_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_899_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_900_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_900_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_900_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_901_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_901_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_901_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_901_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_901_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_902_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_902_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_902_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_903_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_903_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_903_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_903_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_903_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_904_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_904_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_904_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_905_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_905_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_905_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_905_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_905_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_906_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_906_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_906_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_907_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_907_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_907_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_907_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_907_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_908_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_908_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_908_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_909_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_909_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_909_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_909_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_909_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_910_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_910_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_910_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_911_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_911_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_911_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_911_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_911_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_912_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_912_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_912_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_913_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_913_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_913_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_913_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_913_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_914_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_914_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_914_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_915_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_915_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_915_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_915_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_915_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_916_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_916_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_916_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_917_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_917_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_917_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_917_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_917_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_918_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_918_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_918_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_919_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_919_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_919_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_919_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_919_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_920_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_920_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_920_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_921_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_921_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_921_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_921_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_921_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_922_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_922_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_922_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_923_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_923_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_923_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_923_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_923_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_924_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_924_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_924_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_925_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_925_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_925_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_925_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_925_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_926_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_926_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_926_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_927_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_927_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_927_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_927_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_927_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_928_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_928_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_928_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_929_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_929_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_929_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_929_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_929_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_930_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_930_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_930_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_931_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_931_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_931_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_931_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_931_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_932_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_932_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_932_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_933_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_933_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_933_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_933_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_933_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_934_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_934_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_934_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_935_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_935_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_935_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_935_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_935_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_936_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_936_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_936_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_936_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_937_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_937_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_937_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_937_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_937_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_938_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_938_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_938_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_939_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_939_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_939_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_939_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_939_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_940_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_940_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_940_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_941_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_941_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_941_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_941_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_941_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_942_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_942_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_942_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_943_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_943_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_943_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_943_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_943_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_944_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_944_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_944_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_945_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_945_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_945_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_945_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_945_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_946_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_946_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_946_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_947_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_947_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_947_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_947_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_947_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_948_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_948_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_948_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_949_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_949_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_949_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_949_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_949_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_950_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_950_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_950_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_951_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_951_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_951_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_951_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_951_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_952_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_952_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_952_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_953_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_953_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_953_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_953_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_953_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_954_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_954_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_954_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_955_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_955_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_955_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_955_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_955_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_956_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_956_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_956_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_957_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_957_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_957_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_957_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_957_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_958_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_958_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_958_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_959_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_959_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_959_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_959_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_959_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_960_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_960_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_960_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_960_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_961_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_961_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_961_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_961_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_961_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_962_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_962_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_962_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_963_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_963_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_963_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_963_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_963_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_964_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_964_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_964_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_965_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_965_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_965_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_965_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_965_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_966_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_966_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_966_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_967_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_967_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_967_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_967_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_967_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_968_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_968_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_968_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_969_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_969_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_969_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_969_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_969_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_970_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_970_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_970_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_971_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_971_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_971_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_971_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_971_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_972_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_972_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_972_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_973_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_973_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_973_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_973_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_973_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_974_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_974_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_974_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_975_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_975_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_975_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_975_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_975_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_976_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_976_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_976_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_977_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_977_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_977_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_977_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_977_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_978_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_978_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_978_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_979_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_979_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_979_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_979_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_979_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_980_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_980_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_980_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_981_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_981_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_981_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_981_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_981_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_982_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_982_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_982_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_983_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_983_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_983_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_983_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_983_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_984_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_984_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_984_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_985_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_985_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_985_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_985_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_985_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_986_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_986_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_986_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_987_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_987_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_987_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_987_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_987_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_988_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_988_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_988_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_989_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_989_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_989_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_989_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_989_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_990_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_990_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_990_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_991_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_991_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_991_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_991_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_991_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_992_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_992_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_992_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_993_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_993_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_993_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_993_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_993_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_994_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_994_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_994_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_995_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_995_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_995_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_995_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_995_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_996_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_996_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_996_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_997_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_997_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_997_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_997_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_997_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_998_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_998_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_998_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_999_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_999_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_999_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_999_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_999_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_1306 ();
 sky130_fd_sc_hd__decap_3 PHY_1307 ();
 sky130_fd_sc_hd__decap_3 PHY_1308 ();
 sky130_fd_sc_hd__decap_3 PHY_1309 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_1310 ();
 sky130_fd_sc_hd__decap_3 PHY_1311 ();
 sky130_fd_sc_hd__decap_3 PHY_1312 ();
 sky130_fd_sc_hd__decap_3 PHY_1313 ();
 sky130_fd_sc_hd__decap_3 PHY_1314 ();
 sky130_fd_sc_hd__decap_3 PHY_1315 ();
 sky130_fd_sc_hd__decap_3 PHY_1316 ();
 sky130_fd_sc_hd__decap_3 PHY_1317 ();
 sky130_fd_sc_hd__decap_3 PHY_1318 ();
 sky130_fd_sc_hd__decap_3 PHY_1319 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_1320 ();
 sky130_fd_sc_hd__decap_3 PHY_1321 ();
 sky130_fd_sc_hd__decap_3 PHY_1322 ();
 sky130_fd_sc_hd__decap_3 PHY_1323 ();
 sky130_fd_sc_hd__decap_3 PHY_1324 ();
 sky130_fd_sc_hd__decap_3 PHY_1325 ();
 sky130_fd_sc_hd__decap_3 PHY_1326 ();
 sky130_fd_sc_hd__decap_3 PHY_1327 ();
 sky130_fd_sc_hd__decap_3 PHY_1328 ();
 sky130_fd_sc_hd__decap_3 PHY_1329 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_1330 ();
 sky130_fd_sc_hd__decap_3 PHY_1331 ();
 sky130_fd_sc_hd__decap_3 PHY_1332 ();
 sky130_fd_sc_hd__decap_3 PHY_1333 ();
 sky130_fd_sc_hd__decap_3 PHY_1334 ();
 sky130_fd_sc_hd__decap_3 PHY_1335 ();
 sky130_fd_sc_hd__decap_3 PHY_1336 ();
 sky130_fd_sc_hd__decap_3 PHY_1337 ();
 sky130_fd_sc_hd__decap_3 PHY_1338 ();
 sky130_fd_sc_hd__decap_3 PHY_1339 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_1340 ();
 sky130_fd_sc_hd__decap_3 PHY_1341 ();
 sky130_fd_sc_hd__decap_3 PHY_1342 ();
 sky130_fd_sc_hd__decap_3 PHY_1343 ();
 sky130_fd_sc_hd__decap_3 PHY_1344 ();
 sky130_fd_sc_hd__decap_3 PHY_1345 ();
 sky130_fd_sc_hd__decap_3 PHY_1346 ();
 sky130_fd_sc_hd__decap_3 PHY_1347 ();
 sky130_fd_sc_hd__decap_3 PHY_1348 ();
 sky130_fd_sc_hd__decap_3 PHY_1349 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_1350 ();
 sky130_fd_sc_hd__decap_3 PHY_1351 ();
 sky130_fd_sc_hd__decap_3 PHY_1352 ();
 sky130_fd_sc_hd__decap_3 PHY_1353 ();
 sky130_fd_sc_hd__decap_3 PHY_1354 ();
 sky130_fd_sc_hd__decap_3 PHY_1355 ();
 sky130_fd_sc_hd__decap_3 PHY_1356 ();
 sky130_fd_sc_hd__decap_3 PHY_1357 ();
 sky130_fd_sc_hd__decap_3 PHY_1358 ();
 sky130_fd_sc_hd__decap_3 PHY_1359 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_1360 ();
 sky130_fd_sc_hd__decap_3 PHY_1361 ();
 sky130_fd_sc_hd__decap_3 PHY_1362 ();
 sky130_fd_sc_hd__decap_3 PHY_1363 ();
 sky130_fd_sc_hd__decap_3 PHY_1364 ();
 sky130_fd_sc_hd__decap_3 PHY_1365 ();
 sky130_fd_sc_hd__decap_3 PHY_1366 ();
 sky130_fd_sc_hd__decap_3 PHY_1367 ();
 sky130_fd_sc_hd__decap_3 PHY_1368 ();
 sky130_fd_sc_hd__decap_3 PHY_1369 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_1370 ();
 sky130_fd_sc_hd__decap_3 PHY_1371 ();
 sky130_fd_sc_hd__decap_3 PHY_1372 ();
 sky130_fd_sc_hd__decap_3 PHY_1373 ();
 sky130_fd_sc_hd__decap_3 PHY_1374 ();
 sky130_fd_sc_hd__decap_3 PHY_1375 ();
 sky130_fd_sc_hd__decap_3 PHY_1376 ();
 sky130_fd_sc_hd__decap_3 PHY_1377 ();
 sky130_fd_sc_hd__decap_3 PHY_1378 ();
 sky130_fd_sc_hd__decap_3 PHY_1379 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_1380 ();
 sky130_fd_sc_hd__decap_3 PHY_1381 ();
 sky130_fd_sc_hd__decap_3 PHY_1382 ();
 sky130_fd_sc_hd__decap_3 PHY_1383 ();
 sky130_fd_sc_hd__decap_3 PHY_1384 ();
 sky130_fd_sc_hd__decap_3 PHY_1385 ();
 sky130_fd_sc_hd__decap_3 PHY_1386 ();
 sky130_fd_sc_hd__decap_3 PHY_1387 ();
 sky130_fd_sc_hd__decap_3 PHY_1388 ();
 sky130_fd_sc_hd__decap_3 PHY_1389 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_1390 ();
 sky130_fd_sc_hd__decap_3 PHY_1391 ();
 sky130_fd_sc_hd__decap_3 PHY_1392 ();
 sky130_fd_sc_hd__decap_3 PHY_1393 ();
 sky130_fd_sc_hd__decap_3 PHY_1394 ();
 sky130_fd_sc_hd__decap_3 PHY_1395 ();
 sky130_fd_sc_hd__decap_3 PHY_1396 ();
 sky130_fd_sc_hd__decap_3 PHY_1397 ();
 sky130_fd_sc_hd__decap_3 PHY_1398 ();
 sky130_fd_sc_hd__decap_3 PHY_1399 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_1400 ();
 sky130_fd_sc_hd__decap_3 PHY_1401 ();
 sky130_fd_sc_hd__decap_3 PHY_1402 ();
 sky130_fd_sc_hd__decap_3 PHY_1403 ();
 sky130_fd_sc_hd__decap_3 PHY_1404 ();
 sky130_fd_sc_hd__decap_3 PHY_1405 ();
 sky130_fd_sc_hd__decap_3 PHY_1406 ();
 sky130_fd_sc_hd__decap_3 PHY_1407 ();
 sky130_fd_sc_hd__decap_3 PHY_1408 ();
 sky130_fd_sc_hd__decap_3 PHY_1409 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_1410 ();
 sky130_fd_sc_hd__decap_3 PHY_1411 ();
 sky130_fd_sc_hd__decap_3 PHY_1412 ();
 sky130_fd_sc_hd__decap_3 PHY_1413 ();
 sky130_fd_sc_hd__decap_3 PHY_1414 ();
 sky130_fd_sc_hd__decap_3 PHY_1415 ();
 sky130_fd_sc_hd__decap_3 PHY_1416 ();
 sky130_fd_sc_hd__decap_3 PHY_1417 ();
 sky130_fd_sc_hd__decap_3 PHY_1418 ();
 sky130_fd_sc_hd__decap_3 PHY_1419 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_1420 ();
 sky130_fd_sc_hd__decap_3 PHY_1421 ();
 sky130_fd_sc_hd__decap_3 PHY_1422 ();
 sky130_fd_sc_hd__decap_3 PHY_1423 ();
 sky130_fd_sc_hd__decap_3 PHY_1424 ();
 sky130_fd_sc_hd__decap_3 PHY_1425 ();
 sky130_fd_sc_hd__decap_3 PHY_1426 ();
 sky130_fd_sc_hd__decap_3 PHY_1427 ();
 sky130_fd_sc_hd__decap_3 PHY_1428 ();
 sky130_fd_sc_hd__decap_3 PHY_1429 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_1430 ();
 sky130_fd_sc_hd__decap_3 PHY_1431 ();
 sky130_fd_sc_hd__decap_3 PHY_1432 ();
 sky130_fd_sc_hd__decap_3 PHY_1433 ();
 sky130_fd_sc_hd__decap_3 PHY_1434 ();
 sky130_fd_sc_hd__decap_3 PHY_1435 ();
 sky130_fd_sc_hd__decap_3 PHY_1436 ();
 sky130_fd_sc_hd__decap_3 PHY_1437 ();
 sky130_fd_sc_hd__decap_3 PHY_1438 ();
 sky130_fd_sc_hd__decap_3 PHY_1439 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_1440 ();
 sky130_fd_sc_hd__decap_3 PHY_1441 ();
 sky130_fd_sc_hd__decap_3 PHY_1442 ();
 sky130_fd_sc_hd__decap_3 PHY_1443 ();
 sky130_fd_sc_hd__decap_3 PHY_1444 ();
 sky130_fd_sc_hd__decap_3 PHY_1445 ();
 sky130_fd_sc_hd__decap_3 PHY_1446 ();
 sky130_fd_sc_hd__decap_3 PHY_1447 ();
 sky130_fd_sc_hd__decap_3 PHY_1448 ();
 sky130_fd_sc_hd__decap_3 PHY_1449 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_1450 ();
 sky130_fd_sc_hd__decap_3 PHY_1451 ();
 sky130_fd_sc_hd__decap_3 PHY_1452 ();
 sky130_fd_sc_hd__decap_3 PHY_1453 ();
 sky130_fd_sc_hd__decap_3 PHY_1454 ();
 sky130_fd_sc_hd__decap_3 PHY_1455 ();
 sky130_fd_sc_hd__decap_3 PHY_1456 ();
 sky130_fd_sc_hd__decap_3 PHY_1457 ();
 sky130_fd_sc_hd__decap_3 PHY_1458 ();
 sky130_fd_sc_hd__decap_3 PHY_1459 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_1460 ();
 sky130_fd_sc_hd__decap_3 PHY_1461 ();
 sky130_fd_sc_hd__decap_3 PHY_1462 ();
 sky130_fd_sc_hd__decap_3 PHY_1463 ();
 sky130_fd_sc_hd__decap_3 PHY_1464 ();
 sky130_fd_sc_hd__decap_3 PHY_1465 ();
 sky130_fd_sc_hd__decap_3 PHY_1466 ();
 sky130_fd_sc_hd__decap_3 PHY_1467 ();
 sky130_fd_sc_hd__decap_3 PHY_1468 ();
 sky130_fd_sc_hd__decap_3 PHY_1469 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_1470 ();
 sky130_fd_sc_hd__decap_3 PHY_1471 ();
 sky130_fd_sc_hd__decap_3 PHY_1472 ();
 sky130_fd_sc_hd__decap_3 PHY_1473 ();
 sky130_fd_sc_hd__decap_3 PHY_1474 ();
 sky130_fd_sc_hd__decap_3 PHY_1475 ();
 sky130_fd_sc_hd__decap_3 PHY_1476 ();
 sky130_fd_sc_hd__decap_3 PHY_1477 ();
 sky130_fd_sc_hd__decap_3 PHY_1478 ();
 sky130_fd_sc_hd__decap_3 PHY_1479 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_1480 ();
 sky130_fd_sc_hd__decap_3 PHY_1481 ();
 sky130_fd_sc_hd__decap_3 PHY_1482 ();
 sky130_fd_sc_hd__decap_3 PHY_1483 ();
 sky130_fd_sc_hd__decap_3 PHY_1484 ();
 sky130_fd_sc_hd__decap_3 PHY_1485 ();
 sky130_fd_sc_hd__decap_3 PHY_1486 ();
 sky130_fd_sc_hd__decap_3 PHY_1487 ();
 sky130_fd_sc_hd__decap_3 PHY_1488 ();
 sky130_fd_sc_hd__decap_3 PHY_1489 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_1490 ();
 sky130_fd_sc_hd__decap_3 PHY_1491 ();
 sky130_fd_sc_hd__decap_3 PHY_1492 ();
 sky130_fd_sc_hd__decap_3 PHY_1493 ();
 sky130_fd_sc_hd__decap_3 PHY_1494 ();
 sky130_fd_sc_hd__decap_3 PHY_1495 ();
 sky130_fd_sc_hd__decap_3 PHY_1496 ();
 sky130_fd_sc_hd__decap_3 PHY_1497 ();
 sky130_fd_sc_hd__decap_3 PHY_1498 ();
 sky130_fd_sc_hd__decap_3 PHY_1499 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_1500 ();
 sky130_fd_sc_hd__decap_3 PHY_1501 ();
 sky130_fd_sc_hd__decap_3 PHY_1502 ();
 sky130_fd_sc_hd__decap_3 PHY_1503 ();
 sky130_fd_sc_hd__decap_3 PHY_1504 ();
 sky130_fd_sc_hd__decap_3 PHY_1505 ();
 sky130_fd_sc_hd__decap_3 PHY_1506 ();
 sky130_fd_sc_hd__decap_3 PHY_1507 ();
 sky130_fd_sc_hd__decap_3 PHY_1508 ();
 sky130_fd_sc_hd__decap_3 PHY_1509 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_1510 ();
 sky130_fd_sc_hd__decap_3 PHY_1511 ();
 sky130_fd_sc_hd__decap_3 PHY_1512 ();
 sky130_fd_sc_hd__decap_3 PHY_1513 ();
 sky130_fd_sc_hd__decap_3 PHY_1514 ();
 sky130_fd_sc_hd__decap_3 PHY_1515 ();
 sky130_fd_sc_hd__decap_3 PHY_1516 ();
 sky130_fd_sc_hd__decap_3 PHY_1517 ();
 sky130_fd_sc_hd__decap_3 PHY_1518 ();
 sky130_fd_sc_hd__decap_3 PHY_1519 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_1520 ();
 sky130_fd_sc_hd__decap_3 PHY_1521 ();
 sky130_fd_sc_hd__decap_3 PHY_1522 ();
 sky130_fd_sc_hd__decap_3 PHY_1523 ();
 sky130_fd_sc_hd__decap_3 PHY_1524 ();
 sky130_fd_sc_hd__decap_3 PHY_1525 ();
 sky130_fd_sc_hd__decap_3 PHY_1526 ();
 sky130_fd_sc_hd__decap_3 PHY_1527 ();
 sky130_fd_sc_hd__decap_3 PHY_1528 ();
 sky130_fd_sc_hd__decap_3 PHY_1529 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_1530 ();
 sky130_fd_sc_hd__decap_3 PHY_1531 ();
 sky130_fd_sc_hd__decap_3 PHY_1532 ();
 sky130_fd_sc_hd__decap_3 PHY_1533 ();
 sky130_fd_sc_hd__decap_3 PHY_1534 ();
 sky130_fd_sc_hd__decap_3 PHY_1535 ();
 sky130_fd_sc_hd__decap_3 PHY_1536 ();
 sky130_fd_sc_hd__decap_3 PHY_1537 ();
 sky130_fd_sc_hd__decap_3 PHY_1538 ();
 sky130_fd_sc_hd__decap_3 PHY_1539 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_1540 ();
 sky130_fd_sc_hd__decap_3 PHY_1541 ();
 sky130_fd_sc_hd__decap_3 PHY_1542 ();
 sky130_fd_sc_hd__decap_3 PHY_1543 ();
 sky130_fd_sc_hd__decap_3 PHY_1544 ();
 sky130_fd_sc_hd__decap_3 PHY_1545 ();
 sky130_fd_sc_hd__decap_3 PHY_1546 ();
 sky130_fd_sc_hd__decap_3 PHY_1547 ();
 sky130_fd_sc_hd__decap_3 PHY_1548 ();
 sky130_fd_sc_hd__decap_3 PHY_1549 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_1550 ();
 sky130_fd_sc_hd__decap_3 PHY_1551 ();
 sky130_fd_sc_hd__decap_3 PHY_1552 ();
 sky130_fd_sc_hd__decap_3 PHY_1553 ();
 sky130_fd_sc_hd__decap_3 PHY_1554 ();
 sky130_fd_sc_hd__decap_3 PHY_1555 ();
 sky130_fd_sc_hd__decap_3 PHY_1556 ();
 sky130_fd_sc_hd__decap_3 PHY_1557 ();
 sky130_fd_sc_hd__decap_3 PHY_1558 ();
 sky130_fd_sc_hd__decap_3 PHY_1559 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_1560 ();
 sky130_fd_sc_hd__decap_3 PHY_1561 ();
 sky130_fd_sc_hd__decap_3 PHY_1562 ();
 sky130_fd_sc_hd__decap_3 PHY_1563 ();
 sky130_fd_sc_hd__decap_3 PHY_1564 ();
 sky130_fd_sc_hd__decap_3 PHY_1565 ();
 sky130_fd_sc_hd__decap_3 PHY_1566 ();
 sky130_fd_sc_hd__decap_3 PHY_1567 ();
 sky130_fd_sc_hd__decap_3 PHY_1568 ();
 sky130_fd_sc_hd__decap_3 PHY_1569 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_1570 ();
 sky130_fd_sc_hd__decap_3 PHY_1571 ();
 sky130_fd_sc_hd__decap_3 PHY_1572 ();
 sky130_fd_sc_hd__decap_3 PHY_1573 ();
 sky130_fd_sc_hd__decap_3 PHY_1574 ();
 sky130_fd_sc_hd__decap_3 PHY_1575 ();
 sky130_fd_sc_hd__decap_3 PHY_1576 ();
 sky130_fd_sc_hd__decap_3 PHY_1577 ();
 sky130_fd_sc_hd__decap_3 PHY_1578 ();
 sky130_fd_sc_hd__decap_3 PHY_1579 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_1580 ();
 sky130_fd_sc_hd__decap_3 PHY_1581 ();
 sky130_fd_sc_hd__decap_3 PHY_1582 ();
 sky130_fd_sc_hd__decap_3 PHY_1583 ();
 sky130_fd_sc_hd__decap_3 PHY_1584 ();
 sky130_fd_sc_hd__decap_3 PHY_1585 ();
 sky130_fd_sc_hd__decap_3 PHY_1586 ();
 sky130_fd_sc_hd__decap_3 PHY_1587 ();
 sky130_fd_sc_hd__decap_3 PHY_1588 ();
 sky130_fd_sc_hd__decap_3 PHY_1589 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_1590 ();
 sky130_fd_sc_hd__decap_3 PHY_1591 ();
 sky130_fd_sc_hd__decap_3 PHY_1592 ();
 sky130_fd_sc_hd__decap_3 PHY_1593 ();
 sky130_fd_sc_hd__decap_3 PHY_1594 ();
 sky130_fd_sc_hd__decap_3 PHY_1595 ();
 sky130_fd_sc_hd__decap_3 PHY_1596 ();
 sky130_fd_sc_hd__decap_3 PHY_1597 ();
 sky130_fd_sc_hd__decap_3 PHY_1598 ();
 sky130_fd_sc_hd__decap_3 PHY_1599 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_1600 ();
 sky130_fd_sc_hd__decap_3 PHY_1601 ();
 sky130_fd_sc_hd__decap_3 PHY_1602 ();
 sky130_fd_sc_hd__decap_3 PHY_1603 ();
 sky130_fd_sc_hd__decap_3 PHY_1604 ();
 sky130_fd_sc_hd__decap_3 PHY_1605 ();
 sky130_fd_sc_hd__decap_3 PHY_1606 ();
 sky130_fd_sc_hd__decap_3 PHY_1607 ();
 sky130_fd_sc_hd__decap_3 PHY_1608 ();
 sky130_fd_sc_hd__decap_3 PHY_1609 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_1610 ();
 sky130_fd_sc_hd__decap_3 PHY_1611 ();
 sky130_fd_sc_hd__decap_3 PHY_1612 ();
 sky130_fd_sc_hd__decap_3 PHY_1613 ();
 sky130_fd_sc_hd__decap_3 PHY_1614 ();
 sky130_fd_sc_hd__decap_3 PHY_1615 ();
 sky130_fd_sc_hd__decap_3 PHY_1616 ();
 sky130_fd_sc_hd__decap_3 PHY_1617 ();
 sky130_fd_sc_hd__decap_3 PHY_1618 ();
 sky130_fd_sc_hd__decap_3 PHY_1619 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_1620 ();
 sky130_fd_sc_hd__decap_3 PHY_1621 ();
 sky130_fd_sc_hd__decap_3 PHY_1622 ();
 sky130_fd_sc_hd__decap_3 PHY_1623 ();
 sky130_fd_sc_hd__decap_3 PHY_1624 ();
 sky130_fd_sc_hd__decap_3 PHY_1625 ();
 sky130_fd_sc_hd__decap_3 PHY_1626 ();
 sky130_fd_sc_hd__decap_3 PHY_1627 ();
 sky130_fd_sc_hd__decap_3 PHY_1628 ();
 sky130_fd_sc_hd__decap_3 PHY_1629 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_1630 ();
 sky130_fd_sc_hd__decap_3 PHY_1631 ();
 sky130_fd_sc_hd__decap_3 PHY_1632 ();
 sky130_fd_sc_hd__decap_3 PHY_1633 ();
 sky130_fd_sc_hd__decap_3 PHY_1634 ();
 sky130_fd_sc_hd__decap_3 PHY_1635 ();
 sky130_fd_sc_hd__decap_3 PHY_1636 ();
 sky130_fd_sc_hd__decap_3 PHY_1637 ();
 sky130_fd_sc_hd__decap_3 PHY_1638 ();
 sky130_fd_sc_hd__decap_3 PHY_1639 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_1640 ();
 sky130_fd_sc_hd__decap_3 PHY_1641 ();
 sky130_fd_sc_hd__decap_3 PHY_1642 ();
 sky130_fd_sc_hd__decap_3 PHY_1643 ();
 sky130_fd_sc_hd__decap_3 PHY_1644 ();
 sky130_fd_sc_hd__decap_3 PHY_1645 ();
 sky130_fd_sc_hd__decap_3 PHY_1646 ();
 sky130_fd_sc_hd__decap_3 PHY_1647 ();
 sky130_fd_sc_hd__decap_3 PHY_1648 ();
 sky130_fd_sc_hd__decap_3 PHY_1649 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_1650 ();
 sky130_fd_sc_hd__decap_3 PHY_1651 ();
 sky130_fd_sc_hd__decap_3 PHY_1652 ();
 sky130_fd_sc_hd__decap_3 PHY_1653 ();
 sky130_fd_sc_hd__decap_3 PHY_1654 ();
 sky130_fd_sc_hd__decap_3 PHY_1655 ();
 sky130_fd_sc_hd__decap_3 PHY_1656 ();
 sky130_fd_sc_hd__decap_3 PHY_1657 ();
 sky130_fd_sc_hd__decap_3 PHY_1658 ();
 sky130_fd_sc_hd__decap_3 PHY_1659 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_1660 ();
 sky130_fd_sc_hd__decap_3 PHY_1661 ();
 sky130_fd_sc_hd__decap_3 PHY_1662 ();
 sky130_fd_sc_hd__decap_3 PHY_1663 ();
 sky130_fd_sc_hd__decap_3 PHY_1664 ();
 sky130_fd_sc_hd__decap_3 PHY_1665 ();
 sky130_fd_sc_hd__decap_3 PHY_1666 ();
 sky130_fd_sc_hd__decap_3 PHY_1667 ();
 sky130_fd_sc_hd__decap_3 PHY_1668 ();
 sky130_fd_sc_hd__decap_3 PHY_1669 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_1670 ();
 sky130_fd_sc_hd__decap_3 PHY_1671 ();
 sky130_fd_sc_hd__decap_3 PHY_1672 ();
 sky130_fd_sc_hd__decap_3 PHY_1673 ();
 sky130_fd_sc_hd__decap_3 PHY_1674 ();
 sky130_fd_sc_hd__decap_3 PHY_1675 ();
 sky130_fd_sc_hd__decap_3 PHY_1676 ();
 sky130_fd_sc_hd__decap_3 PHY_1677 ();
 sky130_fd_sc_hd__decap_3 PHY_1678 ();
 sky130_fd_sc_hd__decap_3 PHY_1679 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_1680 ();
 sky130_fd_sc_hd__decap_3 PHY_1681 ();
 sky130_fd_sc_hd__decap_3 PHY_1682 ();
 sky130_fd_sc_hd__decap_3 PHY_1683 ();
 sky130_fd_sc_hd__decap_3 PHY_1684 ();
 sky130_fd_sc_hd__decap_3 PHY_1685 ();
 sky130_fd_sc_hd__decap_3 PHY_1686 ();
 sky130_fd_sc_hd__decap_3 PHY_1687 ();
 sky130_fd_sc_hd__decap_3 PHY_1688 ();
 sky130_fd_sc_hd__decap_3 PHY_1689 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_1690 ();
 sky130_fd_sc_hd__decap_3 PHY_1691 ();
 sky130_fd_sc_hd__decap_3 PHY_1692 ();
 sky130_fd_sc_hd__decap_3 PHY_1693 ();
 sky130_fd_sc_hd__decap_3 PHY_1694 ();
 sky130_fd_sc_hd__decap_3 PHY_1695 ();
 sky130_fd_sc_hd__decap_3 PHY_1696 ();
 sky130_fd_sc_hd__decap_3 PHY_1697 ();
 sky130_fd_sc_hd__decap_3 PHY_1698 ();
 sky130_fd_sc_hd__decap_3 PHY_1699 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_1700 ();
 sky130_fd_sc_hd__decap_3 PHY_1701 ();
 sky130_fd_sc_hd__decap_3 PHY_1702 ();
 sky130_fd_sc_hd__decap_3 PHY_1703 ();
 sky130_fd_sc_hd__decap_3 PHY_1704 ();
 sky130_fd_sc_hd__decap_3 PHY_1705 ();
 sky130_fd_sc_hd__decap_3 PHY_1706 ();
 sky130_fd_sc_hd__decap_3 PHY_1707 ();
 sky130_fd_sc_hd__decap_3 PHY_1708 ();
 sky130_fd_sc_hd__decap_3 PHY_1709 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_1710 ();
 sky130_fd_sc_hd__decap_3 PHY_1711 ();
 sky130_fd_sc_hd__decap_3 PHY_1712 ();
 sky130_fd_sc_hd__decap_3 PHY_1713 ();
 sky130_fd_sc_hd__decap_3 PHY_1714 ();
 sky130_fd_sc_hd__decap_3 PHY_1715 ();
 sky130_fd_sc_hd__decap_3 PHY_1716 ();
 sky130_fd_sc_hd__decap_3 PHY_1717 ();
 sky130_fd_sc_hd__decap_3 PHY_1718 ();
 sky130_fd_sc_hd__decap_3 PHY_1719 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_1720 ();
 sky130_fd_sc_hd__decap_3 PHY_1721 ();
 sky130_fd_sc_hd__decap_3 PHY_1722 ();
 sky130_fd_sc_hd__decap_3 PHY_1723 ();
 sky130_fd_sc_hd__decap_3 PHY_1724 ();
 sky130_fd_sc_hd__decap_3 PHY_1725 ();
 sky130_fd_sc_hd__decap_3 PHY_1726 ();
 sky130_fd_sc_hd__decap_3 PHY_1727 ();
 sky130_fd_sc_hd__decap_3 PHY_1728 ();
 sky130_fd_sc_hd__decap_3 PHY_1729 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_1730 ();
 sky130_fd_sc_hd__decap_3 PHY_1731 ();
 sky130_fd_sc_hd__decap_3 PHY_1732 ();
 sky130_fd_sc_hd__decap_3 PHY_1733 ();
 sky130_fd_sc_hd__decap_3 PHY_1734 ();
 sky130_fd_sc_hd__decap_3 PHY_1735 ();
 sky130_fd_sc_hd__decap_3 PHY_1736 ();
 sky130_fd_sc_hd__decap_3 PHY_1737 ();
 sky130_fd_sc_hd__decap_3 PHY_1738 ();
 sky130_fd_sc_hd__decap_3 PHY_1739 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_1740 ();
 sky130_fd_sc_hd__decap_3 PHY_1741 ();
 sky130_fd_sc_hd__decap_3 PHY_1742 ();
 sky130_fd_sc_hd__decap_3 PHY_1743 ();
 sky130_fd_sc_hd__decap_3 PHY_1744 ();
 sky130_fd_sc_hd__decap_3 PHY_1745 ();
 sky130_fd_sc_hd__decap_3 PHY_1746 ();
 sky130_fd_sc_hd__decap_3 PHY_1747 ();
 sky130_fd_sc_hd__decap_3 PHY_1748 ();
 sky130_fd_sc_hd__decap_3 PHY_1749 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_1750 ();
 sky130_fd_sc_hd__decap_3 PHY_1751 ();
 sky130_fd_sc_hd__decap_3 PHY_1752 ();
 sky130_fd_sc_hd__decap_3 PHY_1753 ();
 sky130_fd_sc_hd__decap_3 PHY_1754 ();
 sky130_fd_sc_hd__decap_3 PHY_1755 ();
 sky130_fd_sc_hd__decap_3 PHY_1756 ();
 sky130_fd_sc_hd__decap_3 PHY_1757 ();
 sky130_fd_sc_hd__decap_3 PHY_1758 ();
 sky130_fd_sc_hd__decap_3 PHY_1759 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_1760 ();
 sky130_fd_sc_hd__decap_3 PHY_1761 ();
 sky130_fd_sc_hd__decap_3 PHY_1762 ();
 sky130_fd_sc_hd__decap_3 PHY_1763 ();
 sky130_fd_sc_hd__decap_3 PHY_1764 ();
 sky130_fd_sc_hd__decap_3 PHY_1765 ();
 sky130_fd_sc_hd__decap_3 PHY_1766 ();
 sky130_fd_sc_hd__decap_3 PHY_1767 ();
 sky130_fd_sc_hd__decap_3 PHY_1768 ();
 sky130_fd_sc_hd__decap_3 PHY_1769 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_1770 ();
 sky130_fd_sc_hd__decap_3 PHY_1771 ();
 sky130_fd_sc_hd__decap_3 PHY_1772 ();
 sky130_fd_sc_hd__decap_3 PHY_1773 ();
 sky130_fd_sc_hd__decap_3 PHY_1774 ();
 sky130_fd_sc_hd__decap_3 PHY_1775 ();
 sky130_fd_sc_hd__decap_3 PHY_1776 ();
 sky130_fd_sc_hd__decap_3 PHY_1777 ();
 sky130_fd_sc_hd__decap_3 PHY_1778 ();
 sky130_fd_sc_hd__decap_3 PHY_1779 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_1780 ();
 sky130_fd_sc_hd__decap_3 PHY_1781 ();
 sky130_fd_sc_hd__decap_3 PHY_1782 ();
 sky130_fd_sc_hd__decap_3 PHY_1783 ();
 sky130_fd_sc_hd__decap_3 PHY_1784 ();
 sky130_fd_sc_hd__decap_3 PHY_1785 ();
 sky130_fd_sc_hd__decap_3 PHY_1786 ();
 sky130_fd_sc_hd__decap_3 PHY_1787 ();
 sky130_fd_sc_hd__decap_3 PHY_1788 ();
 sky130_fd_sc_hd__decap_3 PHY_1789 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_1790 ();
 sky130_fd_sc_hd__decap_3 PHY_1791 ();
 sky130_fd_sc_hd__decap_3 PHY_1792 ();
 sky130_fd_sc_hd__decap_3 PHY_1793 ();
 sky130_fd_sc_hd__decap_3 PHY_1794 ();
 sky130_fd_sc_hd__decap_3 PHY_1795 ();
 sky130_fd_sc_hd__decap_3 PHY_1796 ();
 sky130_fd_sc_hd__decap_3 PHY_1797 ();
 sky130_fd_sc_hd__decap_3 PHY_1798 ();
 sky130_fd_sc_hd__decap_3 PHY_1799 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_1800 ();
 sky130_fd_sc_hd__decap_3 PHY_1801 ();
 sky130_fd_sc_hd__decap_3 PHY_1802 ();
 sky130_fd_sc_hd__decap_3 PHY_1803 ();
 sky130_fd_sc_hd__decap_3 PHY_1804 ();
 sky130_fd_sc_hd__decap_3 PHY_1805 ();
 sky130_fd_sc_hd__decap_3 PHY_1806 ();
 sky130_fd_sc_hd__decap_3 PHY_1807 ();
 sky130_fd_sc_hd__decap_3 PHY_1808 ();
 sky130_fd_sc_hd__decap_3 PHY_1809 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_1810 ();
 sky130_fd_sc_hd__decap_3 PHY_1811 ();
 sky130_fd_sc_hd__decap_3 PHY_1812 ();
 sky130_fd_sc_hd__decap_3 PHY_1813 ();
 sky130_fd_sc_hd__decap_3 PHY_1814 ();
 sky130_fd_sc_hd__decap_3 PHY_1815 ();
 sky130_fd_sc_hd__decap_3 PHY_1816 ();
 sky130_fd_sc_hd__decap_3 PHY_1817 ();
 sky130_fd_sc_hd__decap_3 PHY_1818 ();
 sky130_fd_sc_hd__decap_3 PHY_1819 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_1820 ();
 sky130_fd_sc_hd__decap_3 PHY_1821 ();
 sky130_fd_sc_hd__decap_3 PHY_1822 ();
 sky130_fd_sc_hd__decap_3 PHY_1823 ();
 sky130_fd_sc_hd__decap_3 PHY_1824 ();
 sky130_fd_sc_hd__decap_3 PHY_1825 ();
 sky130_fd_sc_hd__decap_3 PHY_1826 ();
 sky130_fd_sc_hd__decap_3 PHY_1827 ();
 sky130_fd_sc_hd__decap_3 PHY_1828 ();
 sky130_fd_sc_hd__decap_3 PHY_1829 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_1830 ();
 sky130_fd_sc_hd__decap_3 PHY_1831 ();
 sky130_fd_sc_hd__decap_3 PHY_1832 ();
 sky130_fd_sc_hd__decap_3 PHY_1833 ();
 sky130_fd_sc_hd__decap_3 PHY_1834 ();
 sky130_fd_sc_hd__decap_3 PHY_1835 ();
 sky130_fd_sc_hd__decap_3 PHY_1836 ();
 sky130_fd_sc_hd__decap_3 PHY_1837 ();
 sky130_fd_sc_hd__decap_3 PHY_1838 ();
 sky130_fd_sc_hd__decap_3 PHY_1839 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_1840 ();
 sky130_fd_sc_hd__decap_3 PHY_1841 ();
 sky130_fd_sc_hd__decap_3 PHY_1842 ();
 sky130_fd_sc_hd__decap_3 PHY_1843 ();
 sky130_fd_sc_hd__decap_3 PHY_1844 ();
 sky130_fd_sc_hd__decap_3 PHY_1845 ();
 sky130_fd_sc_hd__decap_3 PHY_1846 ();
 sky130_fd_sc_hd__decap_3 PHY_1847 ();
 sky130_fd_sc_hd__decap_3 PHY_1848 ();
 sky130_fd_sc_hd__decap_3 PHY_1849 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_1850 ();
 sky130_fd_sc_hd__decap_3 PHY_1851 ();
 sky130_fd_sc_hd__decap_3 PHY_1852 ();
 sky130_fd_sc_hd__decap_3 PHY_1853 ();
 sky130_fd_sc_hd__decap_3 PHY_1854 ();
 sky130_fd_sc_hd__decap_3 PHY_1855 ();
 sky130_fd_sc_hd__decap_3 PHY_1856 ();
 sky130_fd_sc_hd__decap_3 PHY_1857 ();
 sky130_fd_sc_hd__decap_3 PHY_1858 ();
 sky130_fd_sc_hd__decap_3 PHY_1859 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_1860 ();
 sky130_fd_sc_hd__decap_3 PHY_1861 ();
 sky130_fd_sc_hd__decap_3 PHY_1862 ();
 sky130_fd_sc_hd__decap_3 PHY_1863 ();
 sky130_fd_sc_hd__decap_3 PHY_1864 ();
 sky130_fd_sc_hd__decap_3 PHY_1865 ();
 sky130_fd_sc_hd__decap_3 PHY_1866 ();
 sky130_fd_sc_hd__decap_3 PHY_1867 ();
 sky130_fd_sc_hd__decap_3 PHY_1868 ();
 sky130_fd_sc_hd__decap_3 PHY_1869 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_1870 ();
 sky130_fd_sc_hd__decap_3 PHY_1871 ();
 sky130_fd_sc_hd__decap_3 PHY_1872 ();
 sky130_fd_sc_hd__decap_3 PHY_1873 ();
 sky130_fd_sc_hd__decap_3 PHY_1874 ();
 sky130_fd_sc_hd__decap_3 PHY_1875 ();
 sky130_fd_sc_hd__decap_3 PHY_1876 ();
 sky130_fd_sc_hd__decap_3 PHY_1877 ();
 sky130_fd_sc_hd__decap_3 PHY_1878 ();
 sky130_fd_sc_hd__decap_3 PHY_1879 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_1880 ();
 sky130_fd_sc_hd__decap_3 PHY_1881 ();
 sky130_fd_sc_hd__decap_3 PHY_1882 ();
 sky130_fd_sc_hd__decap_3 PHY_1883 ();
 sky130_fd_sc_hd__decap_3 PHY_1884 ();
 sky130_fd_sc_hd__decap_3 PHY_1885 ();
 sky130_fd_sc_hd__decap_3 PHY_1886 ();
 sky130_fd_sc_hd__decap_3 PHY_1887 ();
 sky130_fd_sc_hd__decap_3 PHY_1888 ();
 sky130_fd_sc_hd__decap_3 PHY_1889 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_1890 ();
 sky130_fd_sc_hd__decap_3 PHY_1891 ();
 sky130_fd_sc_hd__decap_3 PHY_1892 ();
 sky130_fd_sc_hd__decap_3 PHY_1893 ();
 sky130_fd_sc_hd__decap_3 PHY_1894 ();
 sky130_fd_sc_hd__decap_3 PHY_1895 ();
 sky130_fd_sc_hd__decap_3 PHY_1896 ();
 sky130_fd_sc_hd__decap_3 PHY_1897 ();
 sky130_fd_sc_hd__decap_3 PHY_1898 ();
 sky130_fd_sc_hd__decap_3 PHY_1899 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_1900 ();
 sky130_fd_sc_hd__decap_3 PHY_1901 ();
 sky130_fd_sc_hd__decap_3 PHY_1902 ();
 sky130_fd_sc_hd__decap_3 PHY_1903 ();
 sky130_fd_sc_hd__decap_3 PHY_1904 ();
 sky130_fd_sc_hd__decap_3 PHY_1905 ();
 sky130_fd_sc_hd__decap_3 PHY_1906 ();
 sky130_fd_sc_hd__decap_3 PHY_1907 ();
 sky130_fd_sc_hd__decap_3 PHY_1908 ();
 sky130_fd_sc_hd__decap_3 PHY_1909 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_1910 ();
 sky130_fd_sc_hd__decap_3 PHY_1911 ();
 sky130_fd_sc_hd__decap_3 PHY_1912 ();
 sky130_fd_sc_hd__decap_3 PHY_1913 ();
 sky130_fd_sc_hd__decap_3 PHY_1914 ();
 sky130_fd_sc_hd__decap_3 PHY_1915 ();
 sky130_fd_sc_hd__decap_3 PHY_1916 ();
 sky130_fd_sc_hd__decap_3 PHY_1917 ();
 sky130_fd_sc_hd__decap_3 PHY_1918 ();
 sky130_fd_sc_hd__decap_3 PHY_1919 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_1920 ();
 sky130_fd_sc_hd__decap_3 PHY_1921 ();
 sky130_fd_sc_hd__decap_3 PHY_1922 ();
 sky130_fd_sc_hd__decap_3 PHY_1923 ();
 sky130_fd_sc_hd__decap_3 PHY_1924 ();
 sky130_fd_sc_hd__decap_3 PHY_1925 ();
 sky130_fd_sc_hd__decap_3 PHY_1926 ();
 sky130_fd_sc_hd__decap_3 PHY_1927 ();
 sky130_fd_sc_hd__decap_3 PHY_1928 ();
 sky130_fd_sc_hd__decap_3 PHY_1929 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_1930 ();
 sky130_fd_sc_hd__decap_3 PHY_1931 ();
 sky130_fd_sc_hd__decap_3 PHY_1932 ();
 sky130_fd_sc_hd__decap_3 PHY_1933 ();
 sky130_fd_sc_hd__decap_3 PHY_1934 ();
 sky130_fd_sc_hd__decap_3 PHY_1935 ();
 sky130_fd_sc_hd__decap_3 PHY_1936 ();
 sky130_fd_sc_hd__decap_3 PHY_1937 ();
 sky130_fd_sc_hd__decap_3 PHY_1938 ();
 sky130_fd_sc_hd__decap_3 PHY_1939 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_1940 ();
 sky130_fd_sc_hd__decap_3 PHY_1941 ();
 sky130_fd_sc_hd__decap_3 PHY_1942 ();
 sky130_fd_sc_hd__decap_3 PHY_1943 ();
 sky130_fd_sc_hd__decap_3 PHY_1944 ();
 sky130_fd_sc_hd__decap_3 PHY_1945 ();
 sky130_fd_sc_hd__decap_3 PHY_1946 ();
 sky130_fd_sc_hd__decap_3 PHY_1947 ();
 sky130_fd_sc_hd__decap_3 PHY_1948 ();
 sky130_fd_sc_hd__decap_3 PHY_1949 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_1950 ();
 sky130_fd_sc_hd__decap_3 PHY_1951 ();
 sky130_fd_sc_hd__decap_3 PHY_1952 ();
 sky130_fd_sc_hd__decap_3 PHY_1953 ();
 sky130_fd_sc_hd__decap_3 PHY_1954 ();
 sky130_fd_sc_hd__decap_3 PHY_1955 ();
 sky130_fd_sc_hd__decap_3 PHY_1956 ();
 sky130_fd_sc_hd__decap_3 PHY_1957 ();
 sky130_fd_sc_hd__decap_3 PHY_1958 ();
 sky130_fd_sc_hd__decap_3 PHY_1959 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_1960 ();
 sky130_fd_sc_hd__decap_3 PHY_1961 ();
 sky130_fd_sc_hd__decap_3 PHY_1962 ();
 sky130_fd_sc_hd__decap_3 PHY_1963 ();
 sky130_fd_sc_hd__decap_3 PHY_1964 ();
 sky130_fd_sc_hd__decap_3 PHY_1965 ();
 sky130_fd_sc_hd__decap_3 PHY_1966 ();
 sky130_fd_sc_hd__decap_3 PHY_1967 ();
 sky130_fd_sc_hd__decap_3 PHY_1968 ();
 sky130_fd_sc_hd__decap_3 PHY_1969 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_1970 ();
 sky130_fd_sc_hd__decap_3 PHY_1971 ();
 sky130_fd_sc_hd__decap_3 PHY_1972 ();
 sky130_fd_sc_hd__decap_3 PHY_1973 ();
 sky130_fd_sc_hd__decap_3 PHY_1974 ();
 sky130_fd_sc_hd__decap_3 PHY_1975 ();
 sky130_fd_sc_hd__decap_3 PHY_1976 ();
 sky130_fd_sc_hd__decap_3 PHY_1977 ();
 sky130_fd_sc_hd__decap_3 PHY_1978 ();
 sky130_fd_sc_hd__decap_3 PHY_1979 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_1980 ();
 sky130_fd_sc_hd__decap_3 PHY_1981 ();
 sky130_fd_sc_hd__decap_3 PHY_1982 ();
 sky130_fd_sc_hd__decap_3 PHY_1983 ();
 sky130_fd_sc_hd__decap_3 PHY_1984 ();
 sky130_fd_sc_hd__decap_3 PHY_1985 ();
 sky130_fd_sc_hd__decap_3 PHY_1986 ();
 sky130_fd_sc_hd__decap_3 PHY_1987 ();
 sky130_fd_sc_hd__decap_3 PHY_1988 ();
 sky130_fd_sc_hd__decap_3 PHY_1989 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_1990 ();
 sky130_fd_sc_hd__decap_3 PHY_1991 ();
 sky130_fd_sc_hd__decap_3 PHY_1992 ();
 sky130_fd_sc_hd__decap_3 PHY_1993 ();
 sky130_fd_sc_hd__decap_3 PHY_1994 ();
 sky130_fd_sc_hd__decap_3 PHY_1995 ();
 sky130_fd_sc_hd__decap_3 PHY_1996 ();
 sky130_fd_sc_hd__decap_3 PHY_1997 ();
 sky130_fd_sc_hd__decap_3 PHY_1998 ();
 sky130_fd_sc_hd__decap_3 PHY_1999 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_2000 ();
 sky130_fd_sc_hd__decap_3 PHY_2001 ();
 sky130_fd_sc_hd__decap_3 PHY_2002 ();
 sky130_fd_sc_hd__decap_3 PHY_2003 ();
 sky130_fd_sc_hd__decap_3 PHY_2004 ();
 sky130_fd_sc_hd__decap_3 PHY_2005 ();
 sky130_fd_sc_hd__decap_3 PHY_2006 ();
 sky130_fd_sc_hd__decap_3 PHY_2007 ();
 sky130_fd_sc_hd__decap_3 PHY_2008 ();
 sky130_fd_sc_hd__decap_3 PHY_2009 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_2010 ();
 sky130_fd_sc_hd__decap_3 PHY_2011 ();
 sky130_fd_sc_hd__decap_3 PHY_2012 ();
 sky130_fd_sc_hd__decap_3 PHY_2013 ();
 sky130_fd_sc_hd__decap_3 PHY_2014 ();
 sky130_fd_sc_hd__decap_3 PHY_2015 ();
 sky130_fd_sc_hd__decap_3 PHY_2016 ();
 sky130_fd_sc_hd__decap_3 PHY_2017 ();
 sky130_fd_sc_hd__decap_3 PHY_2018 ();
 sky130_fd_sc_hd__decap_3 PHY_2019 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_2020 ();
 sky130_fd_sc_hd__decap_3 PHY_2021 ();
 sky130_fd_sc_hd__decap_3 PHY_2022 ();
 sky130_fd_sc_hd__decap_3 PHY_2023 ();
 sky130_fd_sc_hd__decap_3 PHY_2024 ();
 sky130_fd_sc_hd__decap_3 PHY_2025 ();
 sky130_fd_sc_hd__decap_3 PHY_2026 ();
 sky130_fd_sc_hd__decap_3 PHY_2027 ();
 sky130_fd_sc_hd__decap_3 PHY_2028 ();
 sky130_fd_sc_hd__decap_3 PHY_2029 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_2030 ();
 sky130_fd_sc_hd__decap_3 PHY_2031 ();
 sky130_fd_sc_hd__decap_3 PHY_2032 ();
 sky130_fd_sc_hd__decap_3 PHY_2033 ();
 sky130_fd_sc_hd__decap_3 PHY_2034 ();
 sky130_fd_sc_hd__decap_3 PHY_2035 ();
 sky130_fd_sc_hd__decap_3 PHY_2036 ();
 sky130_fd_sc_hd__decap_3 PHY_2037 ();
 sky130_fd_sc_hd__decap_3 PHY_2038 ();
 sky130_fd_sc_hd__decap_3 PHY_2039 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_2040 ();
 sky130_fd_sc_hd__decap_3 PHY_2041 ();
 sky130_fd_sc_hd__decap_3 PHY_2042 ();
 sky130_fd_sc_hd__decap_3 PHY_2043 ();
 sky130_fd_sc_hd__decap_3 PHY_2044 ();
 sky130_fd_sc_hd__decap_3 PHY_2045 ();
 sky130_fd_sc_hd__decap_3 PHY_2046 ();
 sky130_fd_sc_hd__decap_3 PHY_2047 ();
 sky130_fd_sc_hd__decap_3 PHY_2048 ();
 sky130_fd_sc_hd__decap_3 PHY_2049 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_2050 ();
 sky130_fd_sc_hd__decap_3 PHY_2051 ();
 sky130_fd_sc_hd__decap_3 PHY_2052 ();
 sky130_fd_sc_hd__decap_3 PHY_2053 ();
 sky130_fd_sc_hd__decap_3 PHY_2054 ();
 sky130_fd_sc_hd__decap_3 PHY_2055 ();
 sky130_fd_sc_hd__decap_3 PHY_2056 ();
 sky130_fd_sc_hd__decap_3 PHY_2057 ();
 sky130_fd_sc_hd__decap_3 PHY_2058 ();
 sky130_fd_sc_hd__decap_3 PHY_2059 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_2060 ();
 sky130_fd_sc_hd__decap_3 PHY_2061 ();
 sky130_fd_sc_hd__decap_3 PHY_2062 ();
 sky130_fd_sc_hd__decap_3 PHY_2063 ();
 sky130_fd_sc_hd__decap_3 PHY_2064 ();
 sky130_fd_sc_hd__decap_3 PHY_2065 ();
 sky130_fd_sc_hd__decap_3 PHY_2066 ();
 sky130_fd_sc_hd__decap_3 PHY_2067 ();
 sky130_fd_sc_hd__decap_3 PHY_2068 ();
 sky130_fd_sc_hd__decap_3 PHY_2069 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_2070 ();
 sky130_fd_sc_hd__decap_3 PHY_2071 ();
 sky130_fd_sc_hd__decap_3 PHY_2072 ();
 sky130_fd_sc_hd__decap_3 PHY_2073 ();
 sky130_fd_sc_hd__decap_3 PHY_2074 ();
 sky130_fd_sc_hd__decap_3 PHY_2075 ();
 sky130_fd_sc_hd__decap_3 PHY_2076 ();
 sky130_fd_sc_hd__decap_3 PHY_2077 ();
 sky130_fd_sc_hd__decap_3 PHY_2078 ();
 sky130_fd_sc_hd__decap_3 PHY_2079 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_2080 ();
 sky130_fd_sc_hd__decap_3 PHY_2081 ();
 sky130_fd_sc_hd__decap_3 PHY_2082 ();
 sky130_fd_sc_hd__decap_3 PHY_2083 ();
 sky130_fd_sc_hd__decap_3 PHY_2084 ();
 sky130_fd_sc_hd__decap_3 PHY_2085 ();
 sky130_fd_sc_hd__decap_3 PHY_2086 ();
 sky130_fd_sc_hd__decap_3 PHY_2087 ();
 sky130_fd_sc_hd__decap_3 PHY_2088 ();
 sky130_fd_sc_hd__decap_3 PHY_2089 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_2090 ();
 sky130_fd_sc_hd__decap_3 PHY_2091 ();
 sky130_fd_sc_hd__decap_3 PHY_2092 ();
 sky130_fd_sc_hd__decap_3 PHY_2093 ();
 sky130_fd_sc_hd__decap_3 PHY_2094 ();
 sky130_fd_sc_hd__decap_3 PHY_2095 ();
 sky130_fd_sc_hd__decap_3 PHY_2096 ();
 sky130_fd_sc_hd__decap_3 PHY_2097 ();
 sky130_fd_sc_hd__decap_3 PHY_2098 ();
 sky130_fd_sc_hd__decap_3 PHY_2099 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_2100 ();
 sky130_fd_sc_hd__decap_3 PHY_2101 ();
 sky130_fd_sc_hd__decap_3 PHY_2102 ();
 sky130_fd_sc_hd__decap_3 PHY_2103 ();
 sky130_fd_sc_hd__decap_3 PHY_2104 ();
 sky130_fd_sc_hd__decap_3 PHY_2105 ();
 sky130_fd_sc_hd__decap_3 PHY_2106 ();
 sky130_fd_sc_hd__decap_3 PHY_2107 ();
 sky130_fd_sc_hd__decap_3 PHY_2108 ();
 sky130_fd_sc_hd__decap_3 PHY_2109 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_2110 ();
 sky130_fd_sc_hd__decap_3 PHY_2111 ();
 sky130_fd_sc_hd__decap_3 PHY_2112 ();
 sky130_fd_sc_hd__decap_3 PHY_2113 ();
 sky130_fd_sc_hd__decap_3 PHY_2114 ();
 sky130_fd_sc_hd__decap_3 PHY_2115 ();
 sky130_fd_sc_hd__decap_3 PHY_2116 ();
 sky130_fd_sc_hd__decap_3 PHY_2117 ();
 sky130_fd_sc_hd__decap_3 PHY_2118 ();
 sky130_fd_sc_hd__decap_3 PHY_2119 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_2120 ();
 sky130_fd_sc_hd__decap_3 PHY_2121 ();
 sky130_fd_sc_hd__decap_3 PHY_2122 ();
 sky130_fd_sc_hd__decap_3 PHY_2123 ();
 sky130_fd_sc_hd__decap_3 PHY_2124 ();
 sky130_fd_sc_hd__decap_3 PHY_2125 ();
 sky130_fd_sc_hd__decap_3 PHY_2126 ();
 sky130_fd_sc_hd__decap_3 PHY_2127 ();
 sky130_fd_sc_hd__decap_3 PHY_2128 ();
 sky130_fd_sc_hd__decap_3 PHY_2129 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_2130 ();
 sky130_fd_sc_hd__decap_3 PHY_2131 ();
 sky130_fd_sc_hd__decap_3 PHY_2132 ();
 sky130_fd_sc_hd__decap_3 PHY_2133 ();
 sky130_fd_sc_hd__decap_3 PHY_2134 ();
 sky130_fd_sc_hd__decap_3 PHY_2135 ();
 sky130_fd_sc_hd__decap_3 PHY_2136 ();
 sky130_fd_sc_hd__decap_3 PHY_2137 ();
 sky130_fd_sc_hd__decap_3 PHY_2138 ();
 sky130_fd_sc_hd__decap_3 PHY_2139 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_2140 ();
 sky130_fd_sc_hd__decap_3 PHY_2141 ();
 sky130_fd_sc_hd__decap_3 PHY_2142 ();
 sky130_fd_sc_hd__decap_3 PHY_2143 ();
 sky130_fd_sc_hd__decap_3 PHY_2144 ();
 sky130_fd_sc_hd__decap_3 PHY_2145 ();
 sky130_fd_sc_hd__decap_3 PHY_2146 ();
 sky130_fd_sc_hd__decap_3 PHY_2147 ();
 sky130_fd_sc_hd__decap_3 PHY_2148 ();
 sky130_fd_sc_hd__decap_3 PHY_2149 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_2150 ();
 sky130_fd_sc_hd__decap_3 PHY_2151 ();
 sky130_fd_sc_hd__decap_3 PHY_2152 ();
 sky130_fd_sc_hd__decap_3 PHY_2153 ();
 sky130_fd_sc_hd__decap_3 PHY_2154 ();
 sky130_fd_sc_hd__decap_3 PHY_2155 ();
 sky130_fd_sc_hd__decap_3 PHY_2156 ();
 sky130_fd_sc_hd__decap_3 PHY_2157 ();
 sky130_fd_sc_hd__decap_3 PHY_2158 ();
 sky130_fd_sc_hd__decap_3 PHY_2159 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_2160 ();
 sky130_fd_sc_hd__decap_3 PHY_2161 ();
 sky130_fd_sc_hd__decap_3 PHY_2162 ();
 sky130_fd_sc_hd__decap_3 PHY_2163 ();
 sky130_fd_sc_hd__decap_3 PHY_2164 ();
 sky130_fd_sc_hd__decap_3 PHY_2165 ();
 sky130_fd_sc_hd__decap_3 PHY_2166 ();
 sky130_fd_sc_hd__decap_3 PHY_2167 ();
 sky130_fd_sc_hd__decap_3 PHY_2168 ();
 sky130_fd_sc_hd__decap_3 PHY_2169 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_2170 ();
 sky130_fd_sc_hd__decap_3 PHY_2171 ();
 sky130_fd_sc_hd__decap_3 PHY_2172 ();
 sky130_fd_sc_hd__decap_3 PHY_2173 ();
 sky130_fd_sc_hd__decap_3 PHY_2174 ();
 sky130_fd_sc_hd__decap_3 PHY_2175 ();
 sky130_fd_sc_hd__decap_3 PHY_2176 ();
 sky130_fd_sc_hd__decap_3 PHY_2177 ();
 sky130_fd_sc_hd__decap_3 PHY_2178 ();
 sky130_fd_sc_hd__decap_3 PHY_2179 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_2180 ();
 sky130_fd_sc_hd__decap_3 PHY_2181 ();
 sky130_fd_sc_hd__decap_3 PHY_2182 ();
 sky130_fd_sc_hd__decap_3 PHY_2183 ();
 sky130_fd_sc_hd__decap_3 PHY_2184 ();
 sky130_fd_sc_hd__decap_3 PHY_2185 ();
 sky130_fd_sc_hd__decap_3 PHY_2186 ();
 sky130_fd_sc_hd__decap_3 PHY_2187 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__inv_2 _325_ (.A(\Clock_part1.min_tens[3] ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(\Clock_part1.sec_div[8] ),
    .Y(_169_));
 sky130_fd_sc_hd__inv_2 _327_ (.A(\Clock_part1.sec_div[10] ),
    .Y(_170_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(net21),
    .Y(_066_));
 sky130_fd_sc_hd__nand2b_4 _329_ (.A_N(\Clock_part1.dig_cnt[0] ),
    .B(\Clock_part1.dig_cnt[1] ),
    .Y(net5));
 sky130_fd_sc_hd__nand2b_2 _330_ (.A_N(\Clock_part1.dig_cnt[1] ),
    .B(\Clock_part1.dig_cnt[0] ),
    .Y(net4));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(\Clock_part1.scan ),
    .B(\Clock_part1.dig_cnt[0] ),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_8 _332_ (.A(\Clock_part1.dig_cnt[1] ),
    .B(\Clock_part1.dig_cnt[0] ),
    .Y(net6));
 sky130_fd_sc_hd__xnor2_1 _333_ (.A(\Clock_part1.dig_cnt[1] ),
    .B(_171_),
    .Y(_167_));
 sky130_fd_sc_hd__or2_1 _334_ (.A(\Clock_part1.scan ),
    .B(\Clock_part1.dig_cnt[0] ),
    .X(_172_));
 sky130_fd_sc_hd__and2_1 _335_ (.A(_171_),
    .B(_172_),
    .X(_166_));
 sky130_fd_sc_hd__nor3b_2 _336_ (.A(\Clock_part1.min_ones[2] ),
    .B(\Clock_part1.min_ones[1] ),
    .C_N(\Clock_part1.min_ones[3] ),
    .Y(_173_));
 sky130_fd_sc_hd__and4b_1 _337_ (.A_N(\Clock_part1.sec_ones[2] ),
    .B(\Clock_part1.sec_ones[0] ),
    .C(\Clock_part1.sec_ones[3] ),
    .D(\Clock_part1.sec ),
    .X(_174_));
 sky130_fd_sc_hd__and2b_2 _338_ (.A_N(\Clock_part1.sec_ones[1] ),
    .B(_174_),
    .X(_175_));
 sky130_fd_sc_hd__and3b_1 _339_ (.A_N(\Clock_part1.sec_ones[1] ),
    .B(_174_),
    .C(\Clock_part1.sec_tens[0] ),
    .X(_176_));
 sky130_fd_sc_hd__and4bb_1 _340_ (.A_N(\Clock_part1.sec_tens[3] ),
    .B_N(\Clock_part1.sec_tens[1] ),
    .C(_176_),
    .D(\Clock_part1.sec_tens[2] ),
    .X(_177_));
 sky130_fd_sc_hd__and4bb_1 _341_ (.A_N(\Clock_part1.sec_tens[3] ),
    .B_N(\Clock_part1.sec_tens[1] ),
    .C(\Clock_part1.sec_tens[0] ),
    .D(\Clock_part1.sec_tens[2] ),
    .X(_178_));
 sky130_fd_sc_hd__and4b_2 _342_ (.A_N(\Clock_part1.sec_ones[1] ),
    .B(_174_),
    .C(_178_),
    .D(\Clock_part1.min_ones[0] ),
    .X(_179_));
 sky130_fd_sc_hd__and2_1 _343_ (.A(_173_),
    .B(_179_),
    .X(_180_));
 sky130_fd_sc_hd__and3_2 _344_ (.A(\Clock_part1.min_tens[0] ),
    .B(_173_),
    .C(_179_),
    .X(_181_));
 sky130_fd_sc_hd__and4_2 _345_ (.A(\Clock_part1.min_tens[1] ),
    .B(\Clock_part1.min_tens[0] ),
    .C(_173_),
    .D(_179_),
    .X(_182_));
 sky130_fd_sc_hd__nand2_1 _346_ (.A(\Clock_part1.min_tens[2] ),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__and3_1 _347_ (.A(_168_),
    .B(\Clock_part1.min_tens[2] ),
    .C(_182_),
    .X(_184_));
 sky130_fd_sc_hd__a21o_1 _348_ (.A1(\Clock_part1.min_tens[3] ),
    .A2(_183_),
    .B1(_184_),
    .X(_165_));
 sky130_fd_sc_hd__a31oi_4 _349_ (.A1(_168_),
    .A2(\Clock_part1.min_tens[2] ),
    .A3(_181_),
    .B1(_182_),
    .Y(_185_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(_182_),
    .A1(_185_),
    .S(\Clock_part1.min_tens[2] ),
    .X(_164_));
 sky130_fd_sc_hd__o21a_1 _351_ (.A1(\Clock_part1.min_tens[1] ),
    .A2(_181_),
    .B1(_185_),
    .X(_163_));
 sky130_fd_sc_hd__nor2_1 _352_ (.A(\Clock_part1.min_tens[0] ),
    .B(_180_),
    .Y(_186_));
 sky130_fd_sc_hd__nor2_1 _353_ (.A(_181_),
    .B(_186_),
    .Y(_162_));
 sky130_fd_sc_hd__a31oi_1 _354_ (.A1(\Clock_part1.min_ones[2] ),
    .A2(\Clock_part1.min_ones[1] ),
    .A3(_179_),
    .B1(\Clock_part1.min_ones[3] ),
    .Y(_187_));
 sky130_fd_sc_hd__and2_1 _355_ (.A(\Clock_part1.min_ones[1] ),
    .B(_179_),
    .X(_188_));
 sky130_fd_sc_hd__a31o_1 _356_ (.A1(\Clock_part1.min_ones[3] ),
    .A2(\Clock_part1.min_ones[2] ),
    .A3(_188_),
    .B1(_187_),
    .X(_189_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_180_),
    .B(_189_),
    .Y(_161_));
 sky130_fd_sc_hd__xor2_1 _358_ (.A(\Clock_part1.min_ones[2] ),
    .B(_188_),
    .X(_160_));
 sky130_fd_sc_hd__nor2_1 _359_ (.A(\Clock_part1.min_ones[1] ),
    .B(_179_),
    .Y(_190_));
 sky130_fd_sc_hd__nor3_1 _360_ (.A(_173_),
    .B(_188_),
    .C(_190_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _361_ (.A(\Clock_part1.min_ones[0] ),
    .B(_177_),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _362_ (.A(_179_),
    .B(_191_),
    .Y(_158_));
 sky130_fd_sc_hd__and2_1 _363_ (.A(\Clock_part1.sec_tens[1] ),
    .B(_176_),
    .X(_192_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(\Clock_part1.sec_tens[2] ),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__xnor2_1 _365_ (.A(\Clock_part1.sec_tens[3] ),
    .B(_193_),
    .Y(_157_));
 sky130_fd_sc_hd__xnor2_1 _366_ (.A(\Clock_part1.sec_tens[2] ),
    .B(_192_),
    .Y(_194_));
 sky130_fd_sc_hd__nor2_1 _367_ (.A(_177_),
    .B(_194_),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_1 _368_ (.A(\Clock_part1.sec_tens[1] ),
    .B(_176_),
    .Y(_195_));
 sky130_fd_sc_hd__nor3_1 _369_ (.A(_177_),
    .B(_192_),
    .C(_195_),
    .Y(_155_));
 sky130_fd_sc_hd__xor2_1 _370_ (.A(\Clock_part1.sec_tens[0] ),
    .B(_175_),
    .X(_154_));
 sky130_fd_sc_hd__and3_2 _371_ (.A(\Clock_part1.sec ),
    .B(\Clock_part1.sec_ones[1] ),
    .C(\Clock_part1.sec_ones[0] ),
    .X(_196_));
 sky130_fd_sc_hd__a21oi_1 _372_ (.A1(\Clock_part1.sec_ones[2] ),
    .A2(_196_),
    .B1(\Clock_part1.sec_ones[3] ),
    .Y(_197_));
 sky130_fd_sc_hd__a311oi_4 _373_ (.A1(\Clock_part1.sec_ones[3] ),
    .A2(\Clock_part1.sec_ones[2] ),
    .A3(_196_),
    .B1(_197_),
    .C1(_175_),
    .Y(_153_));
 sky130_fd_sc_hd__xor2_1 _374_ (.A(\Clock_part1.sec_ones[2] ),
    .B(_196_),
    .X(_152_));
 sky130_fd_sc_hd__a21oi_1 _375_ (.A1(\Clock_part1.sec ),
    .A2(\Clock_part1.sec_ones[0] ),
    .B1(\Clock_part1.sec_ones[1] ),
    .Y(_198_));
 sky130_fd_sc_hd__nor3_1 _376_ (.A(_174_),
    .B(_196_),
    .C(_198_),
    .Y(_151_));
 sky130_fd_sc_hd__xor2_1 _377_ (.A(\Clock_part1.sec ),
    .B(\Clock_part1.sec_ones[0] ),
    .X(_150_));
 sky130_fd_sc_hd__or4_1 _378_ (.A(\Clock_part1.scan_div[21] ),
    .B(\Clock_part1.scan_div[20] ),
    .C(\Clock_part1.scan_div[23] ),
    .D(\Clock_part1.scan_div[22] ),
    .X(_199_));
 sky130_fd_sc_hd__or4_4 _379_ (.A(\Clock_part1.scan_div[29] ),
    .B(\Clock_part1.scan_div[28] ),
    .C(\Clock_part1.scan_div[31] ),
    .D(\Clock_part1.scan_div[30] ),
    .X(_200_));
 sky130_fd_sc_hd__or4_1 _380_ (.A(\Clock_part1.scan_div[16] ),
    .B(\Clock_part1.scan_div[19] ),
    .C(\Clock_part1.scan_div[24] ),
    .D(\Clock_part1.scan_div[27] ),
    .X(_201_));
 sky130_fd_sc_hd__or4_1 _381_ (.A(\Clock_part1.scan_div[25] ),
    .B(\Clock_part1.scan_div[26] ),
    .C(_200_),
    .D(_201_),
    .X(_202_));
 sky130_fd_sc_hd__or4_1 _382_ (.A(\Clock_part1.scan_div[17] ),
    .B(\Clock_part1.scan_div[18] ),
    .C(_199_),
    .D(_202_),
    .X(_203_));
 sky130_fd_sc_hd__or4b_4 _383_ (.A(\Clock_part1.scan_div[5] ),
    .B(\Clock_part1.scan_div[7] ),
    .C(\Clock_part1.scan_div[6] ),
    .D_N(\Clock_part1.scan_div[4] ),
    .X(_204_));
 sky130_fd_sc_hd__nor2_1 _384_ (.A(\Clock_part1.scan_div[1] ),
    .B(\Clock_part1.scan_div[0] ),
    .Y(_205_));
 sky130_fd_sc_hd__or4bb_1 _385_ (.A(_204_),
    .B(\Clock_part1.scan_div[3] ),
    .C_N(\Clock_part1.scan_div[2] ),
    .D_N(_205_),
    .X(_206_));
 sky130_fd_sc_hd__or4_1 _386_ (.A(\Clock_part1.scan_div[13] ),
    .B(\Clock_part1.scan_div[12] ),
    .C(\Clock_part1.scan_div[15] ),
    .D(\Clock_part1.scan_div[14] ),
    .X(_207_));
 sky130_fd_sc_hd__or4_2 _387_ (.A(\Clock_part1.scan_div[9] ),
    .B(\Clock_part1.scan_div[8] ),
    .C(\Clock_part1.scan_div[11] ),
    .D(\Clock_part1.scan_div[10] ),
    .X(_208_));
 sky130_fd_sc_hd__or4_4 _388_ (.A(_203_),
    .B(_206_),
    .C(_207_),
    .D(_208_),
    .X(_209_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(_209_),
    .Y(_000_));
 sky130_fd_sc_hd__or4_1 _390_ (.A(\Clock_part1.sec_div[21] ),
    .B(\Clock_part1.sec_div[20] ),
    .C(\Clock_part1.sec_div[23] ),
    .D(\Clock_part1.sec_div[22] ),
    .X(_210_));
 sky130_fd_sc_hd__or4_1 _391_ (.A(\Clock_part1.sec_div[17] ),
    .B(\Clock_part1.sec_div[16] ),
    .C(\Clock_part1.sec_div[19] ),
    .D(\Clock_part1.sec_div[18] ),
    .X(_211_));
 sky130_fd_sc_hd__or4_4 _392_ (.A(\Clock_part1.sec_div[25] ),
    .B(\Clock_part1.sec_div[24] ),
    .C(\Clock_part1.sec_div[27] ),
    .D(\Clock_part1.sec_div[26] ),
    .X(_212_));
 sky130_fd_sc_hd__or4_4 _393_ (.A(\Clock_part1.sec_div[29] ),
    .B(\Clock_part1.sec_div[28] ),
    .C(\Clock_part1.sec_div[31] ),
    .D(\Clock_part1.sec_div[30] ),
    .X(_213_));
 sky130_fd_sc_hd__or3_2 _394_ (.A(_210_),
    .B(_211_),
    .C(_213_),
    .X(_214_));
 sky130_fd_sc_hd__or4_4 _395_ (.A(\Clock_part1.sec_div[1] ),
    .B(\Clock_part1.sec_div[0] ),
    .C(\Clock_part1.sec_div[3] ),
    .D(\Clock_part1.sec_div[2] ),
    .X(_215_));
 sky130_fd_sc_hd__nand2_1 _396_ (.A(\Clock_part1.sec_div[6] ),
    .B(\Clock_part1.sec_div[7] ),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_2 _397_ (.A(\Clock_part1.sec_div[8] ),
    .B(\Clock_part1.sec_div[9] ),
    .Y(_217_));
 sky130_fd_sc_hd__or3_1 _398_ (.A(_215_),
    .B(_216_),
    .C(_217_),
    .X(_218_));
 sky130_fd_sc_hd__or4_1 _399_ (.A(\Clock_part1.sec_div[13] ),
    .B(\Clock_part1.sec_div[12] ),
    .C(\Clock_part1.sec_div[15] ),
    .D(\Clock_part1.sec_div[14] ),
    .X(_219_));
 sky130_fd_sc_hd__nand2_1 _400_ (.A(\Clock_part1.sec_div[4] ),
    .B(\Clock_part1.sec_div[10] ),
    .Y(_220_));
 sky130_fd_sc_hd__or4_1 _401_ (.A(\Clock_part1.sec_div[5] ),
    .B(\Clock_part1.sec_div[11] ),
    .C(_219_),
    .D(_220_),
    .X(_221_));
 sky130_fd_sc_hd__or4_4 _402_ (.A(_212_),
    .B(_214_),
    .C(_218_),
    .D(_221_),
    .X(_222_));
 sky130_fd_sc_hd__clkinv_2 _403_ (.A(_222_),
    .Y(_033_));
 sky130_fd_sc_hd__and2b_1 _404_ (.A_N(\Clock_part1.sec_div[0] ),
    .B(_222_),
    .X(_034_));
 sky130_fd_sc_hd__xor2_1 _405_ (.A(\Clock_part1.sec_div[1] ),
    .B(\Clock_part1.sec_div[0] ),
    .X(_045_));
 sky130_fd_sc_hd__and3_1 _406_ (.A(\Clock_part1.sec_div[1] ),
    .B(\Clock_part1.sec_div[0] ),
    .C(\Clock_part1.sec_div[2] ),
    .X(_223_));
 sky130_fd_sc_hd__a21oi_1 _407_ (.A1(\Clock_part1.sec_div[1] ),
    .A2(\Clock_part1.sec_div[0] ),
    .B1(\Clock_part1.sec_div[2] ),
    .Y(_224_));
 sky130_fd_sc_hd__nor2_1 _408_ (.A(_223_),
    .B(_224_),
    .Y(_056_));
 sky130_fd_sc_hd__and4_4 _409_ (.A(\Clock_part1.sec_div[1] ),
    .B(\Clock_part1.sec_div[0] ),
    .C(\Clock_part1.sec_div[3] ),
    .D(\Clock_part1.sec_div[2] ),
    .X(_225_));
 sky130_fd_sc_hd__xor2_1 _410_ (.A(\Clock_part1.sec_div[3] ),
    .B(_223_),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _411_ (.A(\Clock_part1.sec_div[4] ),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__or2_1 _412_ (.A(\Clock_part1.sec_div[4] ),
    .B(_225_),
    .X(_227_));
 sky130_fd_sc_hd__and3_1 _413_ (.A(_222_),
    .B(_226_),
    .C(_227_),
    .X(_060_));
 sky130_fd_sc_hd__xnor2_1 _414_ (.A(\Clock_part1.sec_div[5] ),
    .B(_226_),
    .Y(_061_));
 sky130_fd_sc_hd__a31o_1 _415_ (.A1(\Clock_part1.sec_div[5] ),
    .A2(\Clock_part1.sec_div[4] ),
    .A3(_225_),
    .B1(\Clock_part1.sec_div[6] ),
    .X(_228_));
 sky130_fd_sc_hd__nand4_1 _416_ (.A(\Clock_part1.sec_div[5] ),
    .B(\Clock_part1.sec_div[4] ),
    .C(\Clock_part1.sec_div[6] ),
    .D(_225_),
    .Y(_229_));
 sky130_fd_sc_hd__and3_1 _417_ (.A(_222_),
    .B(_228_),
    .C(_229_),
    .X(_062_));
 sky130_fd_sc_hd__nand2b_1 _418_ (.A_N(\Clock_part1.sec_div[7] ),
    .B(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__and4_1 _419_ (.A(\Clock_part1.sec_div[5] ),
    .B(\Clock_part1.sec_div[4] ),
    .C(\Clock_part1.sec_div[6] ),
    .D(\Clock_part1.sec_div[7] ),
    .X(_231_));
 sky130_fd_sc_hd__nand2_2 _420_ (.A(_225_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__and3_1 _421_ (.A(_222_),
    .B(_230_),
    .C(_232_),
    .X(_063_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_169_),
    .B(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__nor2_1 _423_ (.A(_169_),
    .B(_232_),
    .Y(_234_));
 sky130_fd_sc_hd__o211a_1 _424_ (.A1(_169_),
    .A2(_232_),
    .B1(_233_),
    .C1(_222_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _425_ (.A(\Clock_part1.sec_div[9] ),
    .B(_234_),
    .X(_235_));
 sky130_fd_sc_hd__o211a_1 _426_ (.A1(_217_),
    .A2(_232_),
    .B1(_235_),
    .C1(_222_),
    .X(_065_));
 sky130_fd_sc_hd__o21ai_1 _427_ (.A1(_217_),
    .A2(_232_),
    .B1(_170_),
    .Y(_236_));
 sky130_fd_sc_hd__and3_1 _428_ (.A(\Clock_part1.sec_div[9] ),
    .B(\Clock_part1.sec_div[10] ),
    .C(_234_),
    .X(_237_));
 sky130_fd_sc_hd__o311a_1 _429_ (.A1(_170_),
    .A2(_217_),
    .A3(_232_),
    .B1(_236_),
    .C1(_222_),
    .X(_035_));
 sky130_fd_sc_hd__and4_2 _430_ (.A(\Clock_part1.sec_div[8] ),
    .B(\Clock_part1.sec_div[9] ),
    .C(\Clock_part1.sec_div[11] ),
    .D(\Clock_part1.sec_div[10] ),
    .X(_238_));
 sky130_fd_sc_hd__and3_2 _431_ (.A(_225_),
    .B(_231_),
    .C(_238_),
    .X(_239_));
 sky130_fd_sc_hd__o21ba_1 _432_ (.A1(\Clock_part1.sec_div[11] ),
    .A2(_237_),
    .B1_N(_239_),
    .X(_036_));
 sky130_fd_sc_hd__xor2_1 _433_ (.A(\Clock_part1.sec_div[12] ),
    .B(_239_),
    .X(_037_));
 sky130_fd_sc_hd__and3_1 _434_ (.A(\Clock_part1.sec_div[13] ),
    .B(\Clock_part1.sec_div[12] ),
    .C(_239_),
    .X(_240_));
 sky130_fd_sc_hd__a21o_1 _435_ (.A1(\Clock_part1.sec_div[12] ),
    .A2(_239_),
    .B1(\Clock_part1.sec_div[13] ),
    .X(_241_));
 sky130_fd_sc_hd__and2b_1 _436_ (.A_N(_240_),
    .B(_241_),
    .X(_038_));
 sky130_fd_sc_hd__xor2_1 _437_ (.A(\Clock_part1.sec_div[14] ),
    .B(_240_),
    .X(_039_));
 sky130_fd_sc_hd__a21oi_1 _438_ (.A1(\Clock_part1.sec_div[14] ),
    .A2(_240_),
    .B1(\Clock_part1.sec_div[15] ),
    .Y(_242_));
 sky130_fd_sc_hd__and4_1 _439_ (.A(\Clock_part1.sec_div[13] ),
    .B(\Clock_part1.sec_div[12] ),
    .C(\Clock_part1.sec_div[15] ),
    .D(\Clock_part1.sec_div[14] ),
    .X(_243_));
 sky130_fd_sc_hd__and4_4 _440_ (.A(_225_),
    .B(_231_),
    .C(_238_),
    .D(_243_),
    .X(_244_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(_242_),
    .B(_244_),
    .Y(_040_));
 sky130_fd_sc_hd__xor2_1 _442_ (.A(\Clock_part1.sec_div[16] ),
    .B(_244_),
    .X(_041_));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(\Clock_part1.sec_div[16] ),
    .A2(_244_),
    .B1(\Clock_part1.sec_div[17] ),
    .Y(_245_));
 sky130_fd_sc_hd__and3_1 _444_ (.A(\Clock_part1.sec_div[17] ),
    .B(\Clock_part1.sec_div[16] ),
    .C(_244_),
    .X(_246_));
 sky130_fd_sc_hd__nor2_1 _445_ (.A(_245_),
    .B(_246_),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(\Clock_part1.sec_div[18] ),
    .B(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__and2_1 _447_ (.A(\Clock_part1.sec_div[18] ),
    .B(_246_),
    .X(_248_));
 sky130_fd_sc_hd__nor2_1 _448_ (.A(_247_),
    .B(_248_),
    .Y(_043_));
 sky130_fd_sc_hd__and4_1 _449_ (.A(\Clock_part1.sec_div[17] ),
    .B(\Clock_part1.sec_div[16] ),
    .C(\Clock_part1.sec_div[19] ),
    .D(\Clock_part1.sec_div[18] ),
    .X(_249_));
 sky130_fd_sc_hd__and2_1 _450_ (.A(_244_),
    .B(_249_),
    .X(_250_));
 sky130_fd_sc_hd__o21ba_1 _451_ (.A1(\Clock_part1.sec_div[19] ),
    .A2(_248_),
    .B1_N(_250_),
    .X(_044_));
 sky130_fd_sc_hd__and3_1 _452_ (.A(\Clock_part1.sec_div[20] ),
    .B(_244_),
    .C(_249_),
    .X(_251_));
 sky130_fd_sc_hd__nor2_1 _453_ (.A(\Clock_part1.sec_div[20] ),
    .B(_250_),
    .Y(_252_));
 sky130_fd_sc_hd__nor2_1 _454_ (.A(_251_),
    .B(_252_),
    .Y(_046_));
 sky130_fd_sc_hd__and3_1 _455_ (.A(\Clock_part1.sec_div[21] ),
    .B(\Clock_part1.sec_div[20] ),
    .C(_250_),
    .X(_253_));
 sky130_fd_sc_hd__xor2_1 _456_ (.A(\Clock_part1.sec_div[21] ),
    .B(_251_),
    .X(_047_));
 sky130_fd_sc_hd__xor2_1 _457_ (.A(\Clock_part1.sec_div[22] ),
    .B(_253_),
    .X(_048_));
 sky130_fd_sc_hd__a31o_1 _458_ (.A1(\Clock_part1.sec_div[21] ),
    .A2(\Clock_part1.sec_div[22] ),
    .A3(_251_),
    .B1(\Clock_part1.sec_div[23] ),
    .X(_254_));
 sky130_fd_sc_hd__and4_1 _459_ (.A(\Clock_part1.sec_div[21] ),
    .B(\Clock_part1.sec_div[20] ),
    .C(\Clock_part1.sec_div[23] ),
    .D(\Clock_part1.sec_div[22] ),
    .X(_255_));
 sky130_fd_sc_hd__and3_2 _460_ (.A(_244_),
    .B(_249_),
    .C(_255_),
    .X(_256_));
 sky130_fd_sc_hd__a21boi_1 _461_ (.A1(_250_),
    .A2(_255_),
    .B1_N(_254_),
    .Y(_049_));
 sky130_fd_sc_hd__xor2_1 _462_ (.A(\Clock_part1.sec_div[24] ),
    .B(_256_),
    .X(_050_));
 sky130_fd_sc_hd__and3_1 _463_ (.A(\Clock_part1.sec_div[25] ),
    .B(\Clock_part1.sec_div[24] ),
    .C(_256_),
    .X(_257_));
 sky130_fd_sc_hd__a21o_1 _464_ (.A1(\Clock_part1.sec_div[24] ),
    .A2(_256_),
    .B1(\Clock_part1.sec_div[25] ),
    .X(_258_));
 sky130_fd_sc_hd__and2b_1 _465_ (.A_N(_257_),
    .B(_258_),
    .X(_051_));
 sky130_fd_sc_hd__xor2_1 _466_ (.A(\Clock_part1.sec_div[26] ),
    .B(_257_),
    .X(_052_));
 sky130_fd_sc_hd__and4_1 _467_ (.A(\Clock_part1.sec_div[25] ),
    .B(\Clock_part1.sec_div[24] ),
    .C(\Clock_part1.sec_div[27] ),
    .D(\Clock_part1.sec_div[26] ),
    .X(_259_));
 sky130_fd_sc_hd__and4_2 _468_ (.A(_244_),
    .B(_249_),
    .C(_255_),
    .D(_259_),
    .X(_260_));
 sky130_fd_sc_hd__a41o_1 _469_ (.A1(\Clock_part1.sec_div[25] ),
    .A2(\Clock_part1.sec_div[24] ),
    .A3(\Clock_part1.sec_div[26] ),
    .A4(_256_),
    .B1(\Clock_part1.sec_div[27] ),
    .X(_261_));
 sky130_fd_sc_hd__and2b_1 _470_ (.A_N(_260_),
    .B(_261_),
    .X(_053_));
 sky130_fd_sc_hd__xor2_1 _471_ (.A(\Clock_part1.sec_div[28] ),
    .B(_260_),
    .X(_054_));
 sky130_fd_sc_hd__nand3_1 _472_ (.A(\Clock_part1.sec_div[29] ),
    .B(\Clock_part1.sec_div[28] ),
    .C(_260_),
    .Y(_262_));
 sky130_fd_sc_hd__a21o_1 _473_ (.A1(\Clock_part1.sec_div[28] ),
    .A2(_260_),
    .B1(\Clock_part1.sec_div[29] ),
    .X(_263_));
 sky130_fd_sc_hd__and2_1 _474_ (.A(_262_),
    .B(_263_),
    .X(_055_));
 sky130_fd_sc_hd__and4_1 _475_ (.A(\Clock_part1.sec_div[29] ),
    .B(\Clock_part1.sec_div[28] ),
    .C(\Clock_part1.sec_div[30] ),
    .D(_260_),
    .X(_264_));
 sky130_fd_sc_hd__xnor2_1 _476_ (.A(\Clock_part1.sec_div[30] ),
    .B(_262_),
    .Y(_057_));
 sky130_fd_sc_hd__xor2_1 _477_ (.A(\Clock_part1.sec_div[31] ),
    .B(_264_),
    .X(_058_));
 sky130_fd_sc_hd__and2b_1 _478_ (.A_N(\Clock_part1.scan_div[0] ),
    .B(_209_),
    .X(_001_));
 sky130_fd_sc_hd__and2_1 _479_ (.A(\Clock_part1.scan_div[1] ),
    .B(\Clock_part1.scan_div[0] ),
    .X(_265_));
 sky130_fd_sc_hd__nor2_1 _480_ (.A(_205_),
    .B(_265_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(\Clock_part1.scan_div[2] ),
    .B(_265_),
    .Y(_266_));
 sky130_fd_sc_hd__or2_1 _482_ (.A(\Clock_part1.scan_div[2] ),
    .B(_265_),
    .X(_267_));
 sky130_fd_sc_hd__and3_1 _483_ (.A(_209_),
    .B(_266_),
    .C(_267_),
    .X(_023_));
 sky130_fd_sc_hd__and4_2 _484_ (.A(\Clock_part1.scan_div[1] ),
    .B(\Clock_part1.scan_div[0] ),
    .C(\Clock_part1.scan_div[3] ),
    .D(\Clock_part1.scan_div[2] ),
    .X(_268_));
 sky130_fd_sc_hd__xnor2_1 _485_ (.A(\Clock_part1.scan_div[3] ),
    .B(_266_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(\Clock_part1.scan_div[4] ),
    .B(_268_),
    .Y(_269_));
 sky130_fd_sc_hd__or2_1 _487_ (.A(\Clock_part1.scan_div[4] ),
    .B(_268_),
    .X(_270_));
 sky130_fd_sc_hd__and3_1 _488_ (.A(_209_),
    .B(_269_),
    .C(_270_),
    .X(_027_));
 sky130_fd_sc_hd__xnor2_1 _489_ (.A(\Clock_part1.scan_div[5] ),
    .B(_269_),
    .Y(_028_));
 sky130_fd_sc_hd__and4_1 _490_ (.A(\Clock_part1.scan_div[5] ),
    .B(\Clock_part1.scan_div[4] ),
    .C(\Clock_part1.scan_div[6] ),
    .D(_268_),
    .X(_271_));
 sky130_fd_sc_hd__a31o_1 _491_ (.A1(\Clock_part1.scan_div[5] ),
    .A2(\Clock_part1.scan_div[4] ),
    .A3(_268_),
    .B1(\Clock_part1.scan_div[6] ),
    .X(_272_));
 sky130_fd_sc_hd__and2b_1 _492_ (.A_N(_271_),
    .B(_272_),
    .X(_029_));
 sky130_fd_sc_hd__and4_1 _493_ (.A(\Clock_part1.scan_div[5] ),
    .B(\Clock_part1.scan_div[4] ),
    .C(\Clock_part1.scan_div[7] ),
    .D(\Clock_part1.scan_div[6] ),
    .X(_273_));
 sky130_fd_sc_hd__and2_1 _494_ (.A(_268_),
    .B(_273_),
    .X(_274_));
 sky130_fd_sc_hd__o21ba_1 _495_ (.A1(\Clock_part1.scan_div[7] ),
    .A2(_271_),
    .B1_N(_274_),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _496_ (.A(\Clock_part1.scan_div[8] ),
    .B(_268_),
    .C(_273_),
    .X(_275_));
 sky130_fd_sc_hd__nor2_1 _497_ (.A(\Clock_part1.scan_div[8] ),
    .B(_274_),
    .Y(_276_));
 sky130_fd_sc_hd__nor2_1 _498_ (.A(_275_),
    .B(_276_),
    .Y(_031_));
 sky130_fd_sc_hd__and3_1 _499_ (.A(\Clock_part1.scan_div[9] ),
    .B(\Clock_part1.scan_div[8] ),
    .C(_274_),
    .X(_277_));
 sky130_fd_sc_hd__xor2_1 _500_ (.A(\Clock_part1.scan_div[9] ),
    .B(_275_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _501_ (.A(\Clock_part1.scan_div[10] ),
    .B(_277_),
    .X(_278_));
 sky130_fd_sc_hd__xor2_1 _502_ (.A(\Clock_part1.scan_div[10] ),
    .B(_277_),
    .X(_002_));
 sky130_fd_sc_hd__and4_1 _503_ (.A(\Clock_part1.scan_div[9] ),
    .B(\Clock_part1.scan_div[8] ),
    .C(\Clock_part1.scan_div[11] ),
    .D(\Clock_part1.scan_div[10] ),
    .X(_279_));
 sky130_fd_sc_hd__and3_2 _504_ (.A(_268_),
    .B(_273_),
    .C(_279_),
    .X(_280_));
 sky130_fd_sc_hd__o21ba_1 _505_ (.A1(\Clock_part1.scan_div[11] ),
    .A2(_278_),
    .B1_N(_280_),
    .X(_003_));
 sky130_fd_sc_hd__and2_1 _506_ (.A(\Clock_part1.scan_div[12] ),
    .B(_280_),
    .X(_281_));
 sky130_fd_sc_hd__nor2_1 _507_ (.A(\Clock_part1.scan_div[12] ),
    .B(_280_),
    .Y(_282_));
 sky130_fd_sc_hd__nor2_1 _508_ (.A(_281_),
    .B(_282_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_1 _509_ (.A(\Clock_part1.scan_div[13] ),
    .B(_281_),
    .Y(_283_));
 sky130_fd_sc_hd__and3_1 _510_ (.A(\Clock_part1.scan_div[13] ),
    .B(\Clock_part1.scan_div[12] ),
    .C(_280_),
    .X(_284_));
 sky130_fd_sc_hd__nor2_1 _511_ (.A(_283_),
    .B(_284_),
    .Y(_005_));
 sky130_fd_sc_hd__xor2_1 _512_ (.A(\Clock_part1.scan_div[14] ),
    .B(_284_),
    .X(_006_));
 sky130_fd_sc_hd__a31o_1 _513_ (.A1(\Clock_part1.scan_div[13] ),
    .A2(\Clock_part1.scan_div[14] ),
    .A3(_281_),
    .B1(\Clock_part1.scan_div[15] ),
    .X(_285_));
 sky130_fd_sc_hd__and4_1 _514_ (.A(\Clock_part1.scan_div[13] ),
    .B(\Clock_part1.scan_div[12] ),
    .C(\Clock_part1.scan_div[15] ),
    .D(\Clock_part1.scan_div[14] ),
    .X(_286_));
 sky130_fd_sc_hd__and4_4 _515_ (.A(_268_),
    .B(_273_),
    .C(_279_),
    .D(_286_),
    .X(_287_));
 sky130_fd_sc_hd__a21boi_1 _516_ (.A1(_280_),
    .A2(_286_),
    .B1_N(_285_),
    .Y(_007_));
 sky130_fd_sc_hd__xor2_1 _517_ (.A(\Clock_part1.scan_div[16] ),
    .B(_287_),
    .X(_008_));
 sky130_fd_sc_hd__a21oi_1 _518_ (.A1(\Clock_part1.scan_div[16] ),
    .A2(_287_),
    .B1(\Clock_part1.scan_div[17] ),
    .Y(_288_));
 sky130_fd_sc_hd__and3_1 _519_ (.A(\Clock_part1.scan_div[17] ),
    .B(\Clock_part1.scan_div[16] ),
    .C(_287_),
    .X(_289_));
 sky130_fd_sc_hd__nor2_1 _520_ (.A(_288_),
    .B(_289_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(\Clock_part1.scan_div[18] ),
    .B(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__and2_1 _522_ (.A(\Clock_part1.scan_div[18] ),
    .B(_289_),
    .X(_291_));
 sky130_fd_sc_hd__nor2_1 _523_ (.A(_290_),
    .B(_291_),
    .Y(_010_));
 sky130_fd_sc_hd__and4_1 _524_ (.A(\Clock_part1.scan_div[17] ),
    .B(\Clock_part1.scan_div[16] ),
    .C(\Clock_part1.scan_div[19] ),
    .D(\Clock_part1.scan_div[18] ),
    .X(_292_));
 sky130_fd_sc_hd__and2_1 _525_ (.A(_287_),
    .B(_292_),
    .X(_293_));
 sky130_fd_sc_hd__o21ba_1 _526_ (.A1(\Clock_part1.scan_div[19] ),
    .A2(_291_),
    .B1_N(_293_),
    .X(_011_));
 sky130_fd_sc_hd__and3_1 _527_ (.A(\Clock_part1.scan_div[20] ),
    .B(_287_),
    .C(_292_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(\Clock_part1.scan_div[20] ),
    .B(_293_),
    .Y(_295_));
 sky130_fd_sc_hd__nor2_1 _529_ (.A(_294_),
    .B(_295_),
    .Y(_013_));
 sky130_fd_sc_hd__and3_1 _530_ (.A(\Clock_part1.scan_div[21] ),
    .B(\Clock_part1.scan_div[20] ),
    .C(_293_),
    .X(_296_));
 sky130_fd_sc_hd__xor2_1 _531_ (.A(\Clock_part1.scan_div[21] ),
    .B(_294_),
    .X(_014_));
 sky130_fd_sc_hd__xor2_1 _532_ (.A(\Clock_part1.scan_div[22] ),
    .B(_296_),
    .X(_015_));
 sky130_fd_sc_hd__a31o_1 _533_ (.A1(\Clock_part1.scan_div[21] ),
    .A2(\Clock_part1.scan_div[22] ),
    .A3(_294_),
    .B1(\Clock_part1.scan_div[23] ),
    .X(_297_));
 sky130_fd_sc_hd__and4_1 _534_ (.A(\Clock_part1.scan_div[21] ),
    .B(\Clock_part1.scan_div[20] ),
    .C(\Clock_part1.scan_div[23] ),
    .D(\Clock_part1.scan_div[22] ),
    .X(_298_));
 sky130_fd_sc_hd__and3_2 _535_ (.A(_287_),
    .B(_292_),
    .C(_298_),
    .X(_299_));
 sky130_fd_sc_hd__a21boi_1 _536_ (.A1(_293_),
    .A2(_298_),
    .B1_N(_297_),
    .Y(_016_));
 sky130_fd_sc_hd__nand2_1 _537_ (.A(\Clock_part1.scan_div[24] ),
    .B(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__xor2_1 _538_ (.A(\Clock_part1.scan_div[24] ),
    .B(_299_),
    .X(_017_));
 sky130_fd_sc_hd__and3_1 _539_ (.A(\Clock_part1.scan_div[25] ),
    .B(\Clock_part1.scan_div[24] ),
    .C(_299_),
    .X(_301_));
 sky130_fd_sc_hd__xnor2_1 _540_ (.A(\Clock_part1.scan_div[25] ),
    .B(_300_),
    .Y(_018_));
 sky130_fd_sc_hd__xor2_1 _541_ (.A(\Clock_part1.scan_div[26] ),
    .B(_301_),
    .X(_019_));
 sky130_fd_sc_hd__and4_1 _542_ (.A(\Clock_part1.scan_div[25] ),
    .B(\Clock_part1.scan_div[24] ),
    .C(\Clock_part1.scan_div[27] ),
    .D(\Clock_part1.scan_div[26] ),
    .X(_302_));
 sky130_fd_sc_hd__and4_4 _543_ (.A(_287_),
    .B(_292_),
    .C(_298_),
    .D(_302_),
    .X(_303_));
 sky130_fd_sc_hd__a41o_1 _544_ (.A1(\Clock_part1.scan_div[25] ),
    .A2(\Clock_part1.scan_div[24] ),
    .A3(\Clock_part1.scan_div[26] ),
    .A4(_299_),
    .B1(\Clock_part1.scan_div[27] ),
    .X(_304_));
 sky130_fd_sc_hd__and2b_1 _545_ (.A_N(_303_),
    .B(_304_),
    .X(_020_));
 sky130_fd_sc_hd__xor2_1 _546_ (.A(\Clock_part1.scan_div[28] ),
    .B(_303_),
    .X(_021_));
 sky130_fd_sc_hd__nand3_1 _547_ (.A(\Clock_part1.scan_div[29] ),
    .B(\Clock_part1.scan_div[28] ),
    .C(_303_),
    .Y(_305_));
 sky130_fd_sc_hd__a21o_1 _548_ (.A1(\Clock_part1.scan_div[28] ),
    .A2(_303_),
    .B1(\Clock_part1.scan_div[29] ),
    .X(_306_));
 sky130_fd_sc_hd__and2_1 _549_ (.A(_305_),
    .B(_306_),
    .X(_022_));
 sky130_fd_sc_hd__and4_1 _550_ (.A(\Clock_part1.scan_div[29] ),
    .B(\Clock_part1.scan_div[28] ),
    .C(\Clock_part1.scan_div[30] ),
    .D(_303_),
    .X(_307_));
 sky130_fd_sc_hd__xnor2_1 _551_ (.A(\Clock_part1.scan_div[30] ),
    .B(_305_),
    .Y(_024_));
 sky130_fd_sc_hd__xor2_1 _552_ (.A(\Clock_part1.scan_div[31] ),
    .B(_307_),
    .X(_025_));
 sky130_fd_sc_hd__nor2_2 _553_ (.A(\Clock_part1.dig_cnt[1] ),
    .B(\Clock_part1.dig_cnt[0] ),
    .Y(_308_));
 sky130_fd_sc_hd__inv_4 _554_ (.A(_308_),
    .Y(net2));
 sky130_fd_sc_hd__and3b_1 _555_ (.A_N(\Clock_part1.min_tens[2] ),
    .B(net5),
    .C(net4),
    .X(_309_));
 sky130_fd_sc_hd__o221ai_2 _556_ (.A1(\Clock_part1.min_ones[2] ),
    .A2(net5),
    .B1(net4),
    .B2(\Clock_part1.sec_tens[2] ),
    .C1(net2),
    .Y(_310_));
 sky130_fd_sc_hd__o2bb2a_4 _557_ (.A1_N(\Clock_part1.sec_ones[2] ),
    .A2_N(_308_),
    .B1(_309_),
    .B2(_310_),
    .X(_311_));
 sky130_fd_sc_hd__mux4_2 _558_ (.A0(\Clock_part1.sec_ones[1] ),
    .A1(\Clock_part1.sec_tens[1] ),
    .A2(\Clock_part1.min_ones[1] ),
    .A3(\Clock_part1.min_tens[1] ),
    .S0(\Clock_part1.dig_cnt[0] ),
    .S1(\Clock_part1.dig_cnt[1] ),
    .X(_312_));
 sky130_fd_sc_hd__nand2_1 _559_ (.A(_311_),
    .B(_312_),
    .Y(_313_));
 sky130_fd_sc_hd__nor2_1 _560_ (.A(_311_),
    .B(_312_),
    .Y(_314_));
 sky130_fd_sc_hd__mux4_2 _561_ (.A0(\Clock_part1.sec_ones[0] ),
    .A1(\Clock_part1.sec_tens[0] ),
    .A2(\Clock_part1.min_ones[0] ),
    .A3(\Clock_part1.min_tens[0] ),
    .S0(\Clock_part1.dig_cnt[0] ),
    .S1(\Clock_part1.dig_cnt[1] ),
    .X(_315_));
 sky130_fd_sc_hd__a21oi_2 _562_ (.A1(_312_),
    .A2(_315_),
    .B1(_311_),
    .Y(_316_));
 sky130_fd_sc_hd__o221a_1 _563_ (.A1(\Clock_part1.dig_cnt[1] ),
    .A2(\Clock_part1.sec_tens[3] ),
    .B1(net5),
    .B2(\Clock_part1.min_ones[3] ),
    .C1(net2),
    .X(_317_));
 sky130_fd_sc_hd__or2_1 _564_ (.A(\Clock_part1.min_tens[3] ),
    .B(net6),
    .X(_318_));
 sky130_fd_sc_hd__a22o_4 _565_ (.A1(\Clock_part1.sec_ones[3] ),
    .A2(_308_),
    .B1(_317_),
    .B2(_318_),
    .X(_319_));
 sky130_fd_sc_hd__or3b_1 _566_ (.A(_316_),
    .B(_319_),
    .C_N(_313_),
    .X(net7));
 sky130_fd_sc_hd__or2_1 _567_ (.A(_312_),
    .B(_315_),
    .X(_320_));
 sky130_fd_sc_hd__inv_2 _568_ (.A(_320_),
    .Y(_321_));
 sky130_fd_sc_hd__or3_4 _569_ (.A(_316_),
    .B(_319_),
    .C(_321_),
    .X(net8));
 sky130_fd_sc_hd__nand2b_1 _570_ (.A_N(_312_),
    .B(_311_),
    .Y(_322_));
 sky130_fd_sc_hd__a2bb2o_4 _571_ (.A1_N(_314_),
    .A2_N(_315_),
    .B1(_319_),
    .B2(_322_),
    .X(net9));
 sky130_fd_sc_hd__nand2b_1 _572_ (.A_N(_312_),
    .B(_315_),
    .Y(_323_));
 sky130_fd_sc_hd__a21o_1 _573_ (.A1(_311_),
    .A2(_323_),
    .B1(_319_),
    .X(_324_));
 sky130_fd_sc_hd__a21o_4 _574_ (.A1(_316_),
    .A2(_320_),
    .B1(_324_),
    .X(net10));
 sky130_fd_sc_hd__or3_4 _575_ (.A(_313_),
    .B(_315_),
    .C(_319_),
    .X(net11));
 sky130_fd_sc_hd__or3b_4 _576_ (.A(_319_),
    .B(_321_),
    .C_N(_316_),
    .X(net12));
 sky130_fd_sc_hd__o21bai_4 _577_ (.A1(_311_),
    .A2(_321_),
    .B1_N(_324_),
    .Y(net3));
 sky130_fd_sc_hd__inv_2 _578_ (.A(net19),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _579_ (.A(net21),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(net23),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _581_ (.A(net23),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _582_ (.A(net21),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(net21),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(net21),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _585_ (.A(net13),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _586_ (.A(net13),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _587_ (.A(net17),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _588_ (.A(net17),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _589_ (.A(net13),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _590_ (.A(net14),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _591_ (.A(net13),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _592_ (.A(net14),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _593_ (.A(net15),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _594_ (.A(net15),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _595_ (.A(net15),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _596_ (.A(net15),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _597_ (.A(net19),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _598_ (.A(net19),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _599_ (.A(net19),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _600_ (.A(net18),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _601_ (.A(net18),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _602_ (.A(net19),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _603_ (.A(net19),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _604_ (.A(net18),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _605_ (.A(net21),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _606_ (.A(net23),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _607_ (.A(net23),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _608_ (.A(net23),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _609_ (.A(net21),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _610_ (.A(net21),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _611_ (.A(net21),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _612_ (.A(net21),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _613_ (.A(net15),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _614_ (.A(net17),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _615_ (.A(net17),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _616_ (.A(net15),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _617_ (.A(net13),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _618_ (.A(net14),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _619_ (.A(net13),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _620_ (.A(net13),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _621_ (.A(net13),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _622_ (.A(net14),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _623_ (.A(net14),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _624_ (.A(net13),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _625_ (.A(net15),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _626_ (.A(net16),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _627_ (.A(net16),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _628_ (.A(net16),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _629_ (.A(net18),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _630_ (.A(net15),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _631_ (.A(net15),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _632_ (.A(net17),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _633_ (.A(net17),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _634_ (.A(net17),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _635_ (.A(net13),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _636_ (.A(net14),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _637_ (.A(net18),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _638_ (.A(net16),
    .Y(_127_));
 sky130_fd_sc_hd__inv_2 _639_ (.A(net15),
    .Y(_128_));
 sky130_fd_sc_hd__inv_2 _640_ (.A(net16),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _641_ (.A(net22),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _642_ (.A(net22),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _643_ (.A(net22),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _644_ (.A(net22),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _645_ (.A(net19),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _646_ (.A(net18),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _647_ (.A(net22),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _648_ (.A(net18),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _649_ (.A(net18),
    .Y(_138_));
 sky130_fd_sc_hd__inv_2 _650_ (.A(net20),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _651_ (.A(net20),
    .Y(_140_));
 sky130_fd_sc_hd__inv_2 _652_ (.A(net19),
    .Y(_141_));
 sky130_fd_sc_hd__inv_2 _653_ (.A(net22),
    .Y(_142_));
 sky130_fd_sc_hd__inv_2 _654_ (.A(net19),
    .Y(_143_));
 sky130_fd_sc_hd__inv_2 _655_ (.A(net19),
    .Y(_144_));
 sky130_fd_sc_hd__inv_2 _656_ (.A(net20),
    .Y(_145_));
 sky130_fd_sc_hd__inv_2 _657_ (.A(net23),
    .Y(_146_));
 sky130_fd_sc_hd__inv_2 _658_ (.A(net23),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _659_ (.A(net18),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _660_ (.A(net18),
    .Y(_149_));
 sky130_fd_sc_hd__dfrtp_2 _661_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_150_),
    .RESET_B(_066_),
    .Q(\Clock_part1.sec_ones[0] ));
 sky130_fd_sc_hd__dfrtp_2 _662_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_151_),
    .RESET_B(_067_),
    .Q(\Clock_part1.sec_ones[1] ));
 sky130_fd_sc_hd__dfrtp_4 _663_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_152_),
    .RESET_B(_068_),
    .Q(\Clock_part1.sec_ones[2] ));
 sky130_fd_sc_hd__dfrtp_4 _664_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_153_),
    .RESET_B(_069_),
    .Q(\Clock_part1.sec_ones[3] ));
 sky130_fd_sc_hd__dfrtp_2 _665_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_034_),
    .RESET_B(_070_),
    .Q(\Clock_part1.sec_div[0] ));
 sky130_fd_sc_hd__dfrtp_1 _666_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_045_),
    .RESET_B(_071_),
    .Q(\Clock_part1.sec_div[1] ));
 sky130_fd_sc_hd__dfrtp_1 _667_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_056_),
    .RESET_B(_072_),
    .Q(\Clock_part1.sec_div[2] ));
 sky130_fd_sc_hd__dfrtp_1 _668_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_059_),
    .RESET_B(_073_),
    .Q(\Clock_part1.sec_div[3] ));
 sky130_fd_sc_hd__dfrtp_2 _669_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_060_),
    .RESET_B(_074_),
    .Q(\Clock_part1.sec_div[4] ));
 sky130_fd_sc_hd__dfrtp_2 _670_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_061_),
    .RESET_B(_075_),
    .Q(\Clock_part1.sec_div[5] ));
 sky130_fd_sc_hd__dfrtp_1 _671_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_062_),
    .RESET_B(_076_),
    .Q(\Clock_part1.sec_div[6] ));
 sky130_fd_sc_hd__dfrtp_1 _672_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_063_),
    .RESET_B(_077_),
    .Q(\Clock_part1.sec_div[7] ));
 sky130_fd_sc_hd__dfrtp_1 _673_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_064_),
    .RESET_B(_078_),
    .Q(\Clock_part1.sec_div[8] ));
 sky130_fd_sc_hd__dfrtp_1 _674_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_065_),
    .RESET_B(_079_),
    .Q(\Clock_part1.sec_div[9] ));
 sky130_fd_sc_hd__dfrtp_1 _675_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_035_),
    .RESET_B(_080_),
    .Q(\Clock_part1.sec_div[10] ));
 sky130_fd_sc_hd__dfrtp_1 _676_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_036_),
    .RESET_B(_081_),
    .Q(\Clock_part1.sec_div[11] ));
 sky130_fd_sc_hd__dfrtp_1 _677_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_037_),
    .RESET_B(_082_),
    .Q(\Clock_part1.sec_div[12] ));
 sky130_fd_sc_hd__dfrtp_1 _678_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_038_),
    .RESET_B(_083_),
    .Q(\Clock_part1.sec_div[13] ));
 sky130_fd_sc_hd__dfrtp_1 _679_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_039_),
    .RESET_B(_084_),
    .Q(\Clock_part1.sec_div[14] ));
 sky130_fd_sc_hd__dfrtp_1 _680_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_040_),
    .RESET_B(_085_),
    .Q(\Clock_part1.sec_div[15] ));
 sky130_fd_sc_hd__dfrtp_2 _681_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_041_),
    .RESET_B(_086_),
    .Q(\Clock_part1.sec_div[16] ));
 sky130_fd_sc_hd__dfrtp_1 _682_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_042_),
    .RESET_B(_087_),
    .Q(\Clock_part1.sec_div[17] ));
 sky130_fd_sc_hd__dfrtp_1 _683_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_043_),
    .RESET_B(_088_),
    .Q(\Clock_part1.sec_div[18] ));
 sky130_fd_sc_hd__dfrtp_1 _684_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_044_),
    .RESET_B(_089_),
    .Q(\Clock_part1.sec_div[19] ));
 sky130_fd_sc_hd__dfrtp_1 _685_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_046_),
    .RESET_B(_090_),
    .Q(\Clock_part1.sec_div[20] ));
 sky130_fd_sc_hd__dfrtp_2 _686_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_047_),
    .RESET_B(_091_),
    .Q(\Clock_part1.sec_div[21] ));
 sky130_fd_sc_hd__dfrtp_1 _687_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_048_),
    .RESET_B(_092_),
    .Q(\Clock_part1.sec_div[22] ));
 sky130_fd_sc_hd__dfrtp_1 _688_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_049_),
    .RESET_B(_093_),
    .Q(\Clock_part1.sec_div[23] ));
 sky130_fd_sc_hd__dfrtp_2 _689_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_050_),
    .RESET_B(_094_),
    .Q(\Clock_part1.sec_div[24] ));
 sky130_fd_sc_hd__dfrtp_1 _690_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_051_),
    .RESET_B(_095_),
    .Q(\Clock_part1.sec_div[25] ));
 sky130_fd_sc_hd__dfrtp_1 _691_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_052_),
    .RESET_B(_096_),
    .Q(\Clock_part1.sec_div[26] ));
 sky130_fd_sc_hd__dfrtp_1 _692_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_053_),
    .RESET_B(_097_),
    .Q(\Clock_part1.sec_div[27] ));
 sky130_fd_sc_hd__dfrtp_2 _693_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_054_),
    .RESET_B(_098_),
    .Q(\Clock_part1.sec_div[28] ));
 sky130_fd_sc_hd__dfrtp_1 _694_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_055_),
    .RESET_B(_099_),
    .Q(\Clock_part1.sec_div[29] ));
 sky130_fd_sc_hd__dfrtp_1 _695_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_057_),
    .RESET_B(_100_),
    .Q(\Clock_part1.sec_div[30] ));
 sky130_fd_sc_hd__dfrtp_1 _696_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_058_),
    .RESET_B(_101_),
    .Q(\Clock_part1.sec_div[31] ));
 sky130_fd_sc_hd__dfrtp_1 _697_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_001_),
    .RESET_B(_102_),
    .Q(\Clock_part1.scan_div[0] ));
 sky130_fd_sc_hd__dfrtp_1 _698_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_012_),
    .RESET_B(_103_),
    .Q(\Clock_part1.scan_div[1] ));
 sky130_fd_sc_hd__dfrtp_1 _699_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_023_),
    .RESET_B(_104_),
    .Q(\Clock_part1.scan_div[2] ));
 sky130_fd_sc_hd__dfrtp_1 _700_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_026_),
    .RESET_B(_105_),
    .Q(\Clock_part1.scan_div[3] ));
 sky130_fd_sc_hd__dfrtp_2 _701_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_027_),
    .RESET_B(_106_),
    .Q(\Clock_part1.scan_div[4] ));
 sky130_fd_sc_hd__dfrtp_2 _702_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_028_),
    .RESET_B(_107_),
    .Q(\Clock_part1.scan_div[5] ));
 sky130_fd_sc_hd__dfrtp_1 _703_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_029_),
    .RESET_B(_108_),
    .Q(\Clock_part1.scan_div[6] ));
 sky130_fd_sc_hd__dfrtp_1 _704_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_030_),
    .RESET_B(_109_),
    .Q(\Clock_part1.scan_div[7] ));
 sky130_fd_sc_hd__dfrtp_1 _705_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_031_),
    .RESET_B(_110_),
    .Q(\Clock_part1.scan_div[8] ));
 sky130_fd_sc_hd__dfrtp_1 _706_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_032_),
    .RESET_B(_111_),
    .Q(\Clock_part1.scan_div[9] ));
 sky130_fd_sc_hd__dfrtp_1 _707_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_002_),
    .RESET_B(_112_),
    .Q(\Clock_part1.scan_div[10] ));
 sky130_fd_sc_hd__dfrtp_1 _708_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_003_),
    .RESET_B(_113_),
    .Q(\Clock_part1.scan_div[11] ));
 sky130_fd_sc_hd__dfrtp_1 _709_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_004_),
    .RESET_B(_114_),
    .Q(\Clock_part1.scan_div[12] ));
 sky130_fd_sc_hd__dfrtp_1 _710_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_005_),
    .RESET_B(_115_),
    .Q(\Clock_part1.scan_div[13] ));
 sky130_fd_sc_hd__dfrtp_1 _711_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_006_),
    .RESET_B(_116_),
    .Q(\Clock_part1.scan_div[14] ));
 sky130_fd_sc_hd__dfrtp_1 _712_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_007_),
    .RESET_B(_117_),
    .Q(\Clock_part1.scan_div[15] ));
 sky130_fd_sc_hd__dfrtp_4 _713_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_008_),
    .RESET_B(_118_),
    .Q(\Clock_part1.scan_div[16] ));
 sky130_fd_sc_hd__dfrtp_1 _714_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_009_),
    .RESET_B(_119_),
    .Q(\Clock_part1.scan_div[17] ));
 sky130_fd_sc_hd__dfrtp_1 _715_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_010_),
    .RESET_B(_120_),
    .Q(\Clock_part1.scan_div[18] ));
 sky130_fd_sc_hd__dfrtp_1 _716_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_011_),
    .RESET_B(_121_),
    .Q(\Clock_part1.scan_div[19] ));
 sky130_fd_sc_hd__dfrtp_1 _717_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_013_),
    .RESET_B(_122_),
    .Q(\Clock_part1.scan_div[20] ));
 sky130_fd_sc_hd__dfrtp_1 _718_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_014_),
    .RESET_B(_123_),
    .Q(\Clock_part1.scan_div[21] ));
 sky130_fd_sc_hd__dfrtp_2 _719_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_015_),
    .RESET_B(_124_),
    .Q(\Clock_part1.scan_div[22] ));
 sky130_fd_sc_hd__dfrtp_1 _720_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_016_),
    .RESET_B(_125_),
    .Q(\Clock_part1.scan_div[23] ));
 sky130_fd_sc_hd__dfrtp_4 _721_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_017_),
    .RESET_B(_126_),
    .Q(\Clock_part1.scan_div[24] ));
 sky130_fd_sc_hd__dfrtp_2 _722_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_018_),
    .RESET_B(_127_),
    .Q(\Clock_part1.scan_div[25] ));
 sky130_fd_sc_hd__dfrtp_1 _723_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_019_),
    .RESET_B(_128_),
    .Q(\Clock_part1.scan_div[26] ));
 sky130_fd_sc_hd__dfrtp_1 _724_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_020_),
    .RESET_B(_129_),
    .Q(\Clock_part1.scan_div[27] ));
 sky130_fd_sc_hd__dfrtp_2 _725_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_021_),
    .RESET_B(_130_),
    .Q(\Clock_part1.scan_div[28] ));
 sky130_fd_sc_hd__dfrtp_1 _726_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_022_),
    .RESET_B(_131_),
    .Q(\Clock_part1.scan_div[29] ));
 sky130_fd_sc_hd__dfrtp_1 _727_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_024_),
    .RESET_B(_132_),
    .Q(\Clock_part1.scan_div[30] ));
 sky130_fd_sc_hd__dfrtp_1 _728_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_025_),
    .RESET_B(_133_),
    .Q(\Clock_part1.scan_div[31] ));
 sky130_fd_sc_hd__dfrtp_2 _729_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_033_),
    .RESET_B(_134_),
    .Q(\Clock_part1.sec ));
 sky130_fd_sc_hd__dfrtp_1 _730_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_000_),
    .RESET_B(_135_),
    .Q(\Clock_part1.scan ));
 sky130_fd_sc_hd__dfrtp_4 _731_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_154_),
    .RESET_B(_136_),
    .Q(\Clock_part1.sec_tens[0] ));
 sky130_fd_sc_hd__dfrtp_4 _732_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_155_),
    .RESET_B(_137_),
    .Q(\Clock_part1.sec_tens[1] ));
 sky130_fd_sc_hd__dfrtp_4 _733_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_156_),
    .RESET_B(_138_),
    .Q(\Clock_part1.sec_tens[2] ));
 sky130_fd_sc_hd__dfrtp_4 _734_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_157_),
    .RESET_B(_139_),
    .Q(\Clock_part1.sec_tens[3] ));
 sky130_fd_sc_hd__dfrtp_2 _735_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_158_),
    .RESET_B(_140_),
    .Q(\Clock_part1.min_ones[0] ));
 sky130_fd_sc_hd__dfrtp_2 _736_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_159_),
    .RESET_B(_141_),
    .Q(\Clock_part1.min_ones[1] ));
 sky130_fd_sc_hd__dfrtp_4 _737_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_160_),
    .RESET_B(_142_),
    .Q(\Clock_part1.min_ones[2] ));
 sky130_fd_sc_hd__dfrtp_2 _738_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_161_),
    .RESET_B(_143_),
    .Q(\Clock_part1.min_ones[3] ));
 sky130_fd_sc_hd__dfrtp_1 _739_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_162_),
    .RESET_B(_144_),
    .Q(\Clock_part1.min_tens[0] ));
 sky130_fd_sc_hd__dfrtp_1 _740_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_163_),
    .RESET_B(_145_),
    .Q(\Clock_part1.min_tens[1] ));
 sky130_fd_sc_hd__dfrtp_4 _741_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_164_),
    .RESET_B(_146_),
    .Q(\Clock_part1.min_tens[2] ));
 sky130_fd_sc_hd__dfrtp_1 _742_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_165_),
    .RESET_B(_147_),
    .Q(\Clock_part1.min_tens[3] ));
 sky130_fd_sc_hd__dfrtp_4 _743_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_166_),
    .RESET_B(_148_),
    .Q(\Clock_part1.dig_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _744_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_167_),
    .RESET_B(_149_),
    .Q(\Clock_part1.dig_cnt[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout13 (.A(net24),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net24),
    .X(net14));
 sky130_fd_sc_hd__buf_4 fanout15 (.A(net17),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(net24),
    .X(net17));
 sky130_fd_sc_hd__buf_4 fanout18 (.A(net20),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net24),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout21 (.A(net23),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(net1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__buf_12 output10 (.A(net10),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output11 (.A(net11),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output12 (.A(net12),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_12 output2 (.A(net2),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output3 (.A(net3),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output4 (.A(net4),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output5 (.A(net5),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output6 (.A(net6),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output7 (.A(net7),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output8 (.A(net8),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output9 (.A(net9),
    .X(io_out[6]));
 sky130_fd_sc_hd__conb_1 user_proj_example1_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 user_proj_example1_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 user_proj_example1_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 user_proj_example1_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 user_proj_example1_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 user_proj_example1_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 user_proj_example1_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 user_proj_example1_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 user_proj_example1_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 user_proj_example1_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 user_proj_example1_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 user_proj_example1_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 user_proj_example1_37 (.HI(net37));
 assign io_oeb[0] = net25;
 assign io_oeb[10] = net35;
 assign io_oeb[11] = net36;
 assign io_oeb[1] = net26;
 assign io_oeb[2] = net27;
 assign io_oeb[3] = net28;
 assign io_oeb[4] = net29;
 assign io_oeb[5] = net30;
 assign io_oeb[6] = net31;
 assign io_oeb[7] = net32;
 assign io_oeb[8] = net33;
 assign io_oeb[9] = net34;
 assign io_out[11] = net37;
endmodule


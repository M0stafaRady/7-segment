VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example1
  CLASS BLOCK ;
  FOREIGN user_proj_example1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 76.200 200.000 76.800 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.000 4.000 1375.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END io_in[11]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 447.480 200.000 448.080 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 818.760 200.000 819.360 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1190.040 200.000 1190.640 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1561.320 200.000 1561.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1932.600 200.000 1933.200 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2303.880 200.000 2304.480 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2675.160 200.000 2675.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2868.280 4.000 2868.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2121.640 4.000 2122.240 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 323.720 200.000 324.320 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[11]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 695.000 200.000 695.600 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1066.280 200.000 1066.880 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1437.560 200.000 1438.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1808.840 200.000 1809.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2180.120 200.000 2180.720 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2551.400 200.000 2552.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2922.680 200.000 2923.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2370.520 4.000 2371.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1623.880 4.000 1624.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 199.960 200.000 200.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.120 4.000 1126.720 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END io_out[11]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 571.240 200.000 571.840 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 942.520 200.000 943.120 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1313.800 200.000 1314.400 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1685.080 200.000 1685.680 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2056.360 200.000 2056.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2427.640 200.000 2428.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2798.920 200.000 2799.520 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2619.400 4.000 2620.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1872.760 4.000 1873.360 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.120 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 192.650 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 192.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 2923.680 196.000 2986.725 ;
        RECT 4.000 2922.280 195.600 2923.680 ;
        RECT 4.000 2869.280 196.000 2922.280 ;
        RECT 4.400 2867.880 196.000 2869.280 ;
        RECT 4.000 2799.920 196.000 2867.880 ;
        RECT 4.000 2798.520 195.600 2799.920 ;
        RECT 4.000 2676.160 196.000 2798.520 ;
        RECT 4.000 2674.760 195.600 2676.160 ;
        RECT 4.000 2620.400 196.000 2674.760 ;
        RECT 4.400 2619.000 196.000 2620.400 ;
        RECT 4.000 2552.400 196.000 2619.000 ;
        RECT 4.000 2551.000 195.600 2552.400 ;
        RECT 4.000 2428.640 196.000 2551.000 ;
        RECT 4.000 2427.240 195.600 2428.640 ;
        RECT 4.000 2371.520 196.000 2427.240 ;
        RECT 4.400 2370.120 196.000 2371.520 ;
        RECT 4.000 2304.880 196.000 2370.120 ;
        RECT 4.000 2303.480 195.600 2304.880 ;
        RECT 4.000 2181.120 196.000 2303.480 ;
        RECT 4.000 2179.720 195.600 2181.120 ;
        RECT 4.000 2122.640 196.000 2179.720 ;
        RECT 4.400 2121.240 196.000 2122.640 ;
        RECT 4.000 2057.360 196.000 2121.240 ;
        RECT 4.000 2055.960 195.600 2057.360 ;
        RECT 4.000 1933.600 196.000 2055.960 ;
        RECT 4.000 1932.200 195.600 1933.600 ;
        RECT 4.000 1873.760 196.000 1932.200 ;
        RECT 4.400 1872.360 196.000 1873.760 ;
        RECT 4.000 1809.840 196.000 1872.360 ;
        RECT 4.000 1808.440 195.600 1809.840 ;
        RECT 4.000 1686.080 196.000 1808.440 ;
        RECT 4.000 1684.680 195.600 1686.080 ;
        RECT 4.000 1624.880 196.000 1684.680 ;
        RECT 4.400 1623.480 196.000 1624.880 ;
        RECT 4.000 1562.320 196.000 1623.480 ;
        RECT 4.000 1560.920 195.600 1562.320 ;
        RECT 4.000 1438.560 196.000 1560.920 ;
        RECT 4.000 1437.160 195.600 1438.560 ;
        RECT 4.000 1376.000 196.000 1437.160 ;
        RECT 4.400 1374.600 196.000 1376.000 ;
        RECT 4.000 1314.800 196.000 1374.600 ;
        RECT 4.000 1313.400 195.600 1314.800 ;
        RECT 4.000 1191.040 196.000 1313.400 ;
        RECT 4.000 1189.640 195.600 1191.040 ;
        RECT 4.000 1127.120 196.000 1189.640 ;
        RECT 4.400 1125.720 196.000 1127.120 ;
        RECT 4.000 1067.280 196.000 1125.720 ;
        RECT 4.000 1065.880 195.600 1067.280 ;
        RECT 4.000 943.520 196.000 1065.880 ;
        RECT 4.000 942.120 195.600 943.520 ;
        RECT 4.000 878.240 196.000 942.120 ;
        RECT 4.400 876.840 196.000 878.240 ;
        RECT 4.000 819.760 196.000 876.840 ;
        RECT 4.000 818.360 195.600 819.760 ;
        RECT 4.000 696.000 196.000 818.360 ;
        RECT 4.000 694.600 195.600 696.000 ;
        RECT 4.000 629.360 196.000 694.600 ;
        RECT 4.400 627.960 196.000 629.360 ;
        RECT 4.000 572.240 196.000 627.960 ;
        RECT 4.000 570.840 195.600 572.240 ;
        RECT 4.000 448.480 196.000 570.840 ;
        RECT 4.000 447.080 195.600 448.480 ;
        RECT 4.000 380.480 196.000 447.080 ;
        RECT 4.400 379.080 196.000 380.480 ;
        RECT 4.000 324.720 196.000 379.080 ;
        RECT 4.000 323.320 195.600 324.720 ;
        RECT 4.000 200.960 196.000 323.320 ;
        RECT 4.000 199.560 195.600 200.960 ;
        RECT 4.000 131.600 196.000 199.560 ;
        RECT 4.400 130.200 196.000 131.600 ;
        RECT 4.000 77.200 196.000 130.200 ;
        RECT 4.000 75.800 195.600 77.200 ;
        RECT 4.000 10.715 196.000 75.800 ;
  END
END user_proj_example1
END LIBRARY


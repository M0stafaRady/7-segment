magic
tech sky130A
magscale 1 2
timestamp 1687358410
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 934 2128 38824 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 938 856 38530 597349
rect 938 800 9898 856
rect 10066 800 29862 856
rect 30030 800 38530 856
<< metal3 >>
rect 39200 584536 40000 584656
rect 0 573656 800 573776
rect 39200 559784 40000 559904
rect 39200 535032 40000 535152
rect 0 523880 800 524000
rect 39200 510280 40000 510400
rect 39200 485528 40000 485648
rect 0 474104 800 474224
rect 39200 460776 40000 460896
rect 39200 436024 40000 436144
rect 0 424328 800 424448
rect 39200 411272 40000 411392
rect 39200 386520 40000 386640
rect 0 374552 800 374672
rect 39200 361768 40000 361888
rect 39200 337016 40000 337136
rect 0 324776 800 324896
rect 39200 312264 40000 312384
rect 39200 287512 40000 287632
rect 0 275000 800 275120
rect 39200 262760 40000 262880
rect 39200 238008 40000 238128
rect 0 225224 800 225344
rect 39200 213256 40000 213376
rect 39200 188504 40000 188624
rect 0 175448 800 175568
rect 39200 163752 40000 163872
rect 39200 139000 40000 139120
rect 0 125672 800 125792
rect 39200 114248 40000 114368
rect 39200 89496 40000 89616
rect 0 75896 800 76016
rect 39200 64744 40000 64864
rect 39200 39992 40000 40112
rect 0 26120 800 26240
rect 39200 15240 40000 15360
<< obsm3 >>
rect 800 584736 39200 597345
rect 800 584456 39120 584736
rect 800 573856 39200 584456
rect 880 573576 39200 573856
rect 800 559984 39200 573576
rect 800 559704 39120 559984
rect 800 535232 39200 559704
rect 800 534952 39120 535232
rect 800 524080 39200 534952
rect 880 523800 39200 524080
rect 800 510480 39200 523800
rect 800 510200 39120 510480
rect 800 485728 39200 510200
rect 800 485448 39120 485728
rect 800 474304 39200 485448
rect 880 474024 39200 474304
rect 800 460976 39200 474024
rect 800 460696 39120 460976
rect 800 436224 39200 460696
rect 800 435944 39120 436224
rect 800 424528 39200 435944
rect 880 424248 39200 424528
rect 800 411472 39200 424248
rect 800 411192 39120 411472
rect 800 386720 39200 411192
rect 800 386440 39120 386720
rect 800 374752 39200 386440
rect 880 374472 39200 374752
rect 800 361968 39200 374472
rect 800 361688 39120 361968
rect 800 337216 39200 361688
rect 800 336936 39120 337216
rect 800 324976 39200 336936
rect 880 324696 39200 324976
rect 800 312464 39200 324696
rect 800 312184 39120 312464
rect 800 287712 39200 312184
rect 800 287432 39120 287712
rect 800 275200 39200 287432
rect 880 274920 39200 275200
rect 800 262960 39200 274920
rect 800 262680 39120 262960
rect 800 238208 39200 262680
rect 800 237928 39120 238208
rect 800 225424 39200 237928
rect 880 225144 39200 225424
rect 800 213456 39200 225144
rect 800 213176 39120 213456
rect 800 188704 39200 213176
rect 800 188424 39120 188704
rect 800 175648 39200 188424
rect 880 175368 39200 175648
rect 800 163952 39200 175368
rect 800 163672 39120 163952
rect 800 139200 39200 163672
rect 800 138920 39120 139200
rect 800 125872 39200 138920
rect 880 125592 39200 125872
rect 800 114448 39200 125592
rect 800 114168 39120 114448
rect 800 89696 39200 114168
rect 800 89416 39120 89696
rect 800 76096 39200 89416
rect 880 75816 39200 76096
rect 800 64944 39200 75816
rect 800 64664 39120 64944
rect 800 40192 39200 64664
rect 800 39912 39120 40192
rect 800 26320 39200 39912
rect 880 26040 39200 26320
rect 800 15440 39200 26040
rect 800 15160 39120 15440
rect 800 2143 39200 15160
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< labels >>
rlabel metal3 s 39200 15240 40000 15360 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 275000 800 275120 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 89496 40000 89616 6 io_in[1]
port 4 nsew signal input
rlabel metal3 s 39200 163752 40000 163872 6 io_in[2]
port 5 nsew signal input
rlabel metal3 s 39200 238008 40000 238128 6 io_in[3]
port 6 nsew signal input
rlabel metal3 s 39200 312264 40000 312384 6 io_in[4]
port 7 nsew signal input
rlabel metal3 s 39200 386520 40000 386640 6 io_in[5]
port 8 nsew signal input
rlabel metal3 s 39200 460776 40000 460896 6 io_in[6]
port 9 nsew signal input
rlabel metal3 s 39200 535032 40000 535152 6 io_in[7]
port 10 nsew signal input
rlabel metal3 s 0 573656 800 573776 6 io_in[8]
port 11 nsew signal input
rlabel metal3 s 0 424328 800 424448 6 io_in[9]
port 12 nsew signal input
rlabel metal3 s 39200 64744 40000 64864 6 io_oeb[0]
port 13 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 io_oeb[10]
port 14 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[11]
port 15 nsew signal output
rlabel metal3 s 39200 139000 40000 139120 6 io_oeb[1]
port 16 nsew signal output
rlabel metal3 s 39200 213256 40000 213376 6 io_oeb[2]
port 17 nsew signal output
rlabel metal3 s 39200 287512 40000 287632 6 io_oeb[3]
port 18 nsew signal output
rlabel metal3 s 39200 361768 40000 361888 6 io_oeb[4]
port 19 nsew signal output
rlabel metal3 s 39200 436024 40000 436144 6 io_oeb[5]
port 20 nsew signal output
rlabel metal3 s 39200 510280 40000 510400 6 io_oeb[6]
port 21 nsew signal output
rlabel metal3 s 39200 584536 40000 584656 6 io_oeb[7]
port 22 nsew signal output
rlabel metal3 s 0 474104 800 474224 6 io_oeb[8]
port 23 nsew signal output
rlabel metal3 s 0 324776 800 324896 6 io_oeb[9]
port 24 nsew signal output
rlabel metal3 s 39200 39992 40000 40112 6 io_out[0]
port 25 nsew signal output
rlabel metal3 s 0 225224 800 225344 6 io_out[10]
port 26 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 io_out[11]
port 27 nsew signal output
rlabel metal3 s 39200 114248 40000 114368 6 io_out[1]
port 28 nsew signal output
rlabel metal3 s 39200 188504 40000 188624 6 io_out[2]
port 29 nsew signal output
rlabel metal3 s 39200 262760 40000 262880 6 io_out[3]
port 30 nsew signal output
rlabel metal3 s 39200 337016 40000 337136 6 io_out[4]
port 31 nsew signal output
rlabel metal3 s 39200 411272 40000 411392 6 io_out[5]
port 32 nsew signal output
rlabel metal3 s 39200 485528 40000 485648 6 io_out[6]
port 33 nsew signal output
rlabel metal3 s 39200 559784 40000 559904 6 io_out[7]
port 34 nsew signal output
rlabel metal3 s 0 523880 800 524000 6 io_out[8]
port 35 nsew signal output
rlabel metal3 s 0 374552 800 374672 6 io_out[9]
port 36 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 38 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 39 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 40 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7604106
string GDS_FILE /home/hosni/OpenLane-tutorial/7-segment/openlane/user_proj_example1/runs/23_06_21_07_38/results/signoff/user_proj_example1.magic.gds
string GDS_START 472770
<< end >>


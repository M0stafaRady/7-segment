magic
tech sky130A
magscale 1 2
timestamp 1687356621
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 934 2128 39086 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 938 856 39082 597349
rect 938 800 9898 856
rect 10066 800 29862 856
rect 30030 800 39082 856
<< metal3 >>
rect 39200 586168 40000 586288
rect 0 574472 800 574592
rect 39200 561280 40000 561400
rect 39200 536392 40000 536512
rect 0 524560 800 524680
rect 39200 511504 40000 511624
rect 39200 486616 40000 486736
rect 0 474648 800 474768
rect 39200 461728 40000 461848
rect 39200 436840 40000 436960
rect 0 424736 800 424856
rect 39200 411952 40000 412072
rect 39200 387064 40000 387184
rect 0 374824 800 374944
rect 39200 362176 40000 362296
rect 39200 337288 40000 337408
rect 0 324912 800 325032
rect 39200 312400 40000 312520
rect 39200 287512 40000 287632
rect 0 275000 800 275120
rect 39200 262624 40000 262744
rect 39200 237736 40000 237856
rect 0 225088 800 225208
rect 39200 212848 40000 212968
rect 39200 187960 40000 188080
rect 0 175176 800 175296
rect 39200 163072 40000 163192
rect 39200 138184 40000 138304
rect 0 125264 800 125384
rect 39200 113296 40000 113416
rect 39200 88408 40000 88528
rect 0 75352 800 75472
rect 39200 63520 40000 63640
rect 39200 38632 40000 38752
rect 0 25440 800 25560
rect 39200 13744 40000 13864
<< obsm3 >>
rect 800 586368 39200 597345
rect 800 586088 39120 586368
rect 800 574672 39200 586088
rect 880 574392 39200 574672
rect 800 561480 39200 574392
rect 800 561200 39120 561480
rect 800 536592 39200 561200
rect 800 536312 39120 536592
rect 800 524760 39200 536312
rect 880 524480 39200 524760
rect 800 511704 39200 524480
rect 800 511424 39120 511704
rect 800 486816 39200 511424
rect 800 486536 39120 486816
rect 800 474848 39200 486536
rect 880 474568 39200 474848
rect 800 461928 39200 474568
rect 800 461648 39120 461928
rect 800 437040 39200 461648
rect 800 436760 39120 437040
rect 800 424936 39200 436760
rect 880 424656 39200 424936
rect 800 412152 39200 424656
rect 800 411872 39120 412152
rect 800 387264 39200 411872
rect 800 386984 39120 387264
rect 800 375024 39200 386984
rect 880 374744 39200 375024
rect 800 362376 39200 374744
rect 800 362096 39120 362376
rect 800 337488 39200 362096
rect 800 337208 39120 337488
rect 800 325112 39200 337208
rect 880 324832 39200 325112
rect 800 312600 39200 324832
rect 800 312320 39120 312600
rect 800 287712 39200 312320
rect 800 287432 39120 287712
rect 800 275200 39200 287432
rect 880 274920 39200 275200
rect 800 262824 39200 274920
rect 800 262544 39120 262824
rect 800 237936 39200 262544
rect 800 237656 39120 237936
rect 800 225288 39200 237656
rect 880 225008 39200 225288
rect 800 213048 39200 225008
rect 800 212768 39120 213048
rect 800 188160 39200 212768
rect 800 187880 39120 188160
rect 800 175376 39200 187880
rect 880 175096 39200 175376
rect 800 163272 39200 175096
rect 800 162992 39120 163272
rect 800 138384 39200 162992
rect 800 138104 39120 138384
rect 800 125464 39200 138104
rect 880 125184 39200 125464
rect 800 113496 39200 125184
rect 800 113216 39120 113496
rect 800 88608 39200 113216
rect 800 88328 39120 88608
rect 800 75552 39200 88328
rect 880 75272 39200 75552
rect 800 63720 39200 75272
rect 800 63440 39120 63720
rect 800 38832 39200 63440
rect 800 38552 39120 38832
rect 800 25640 39200 38552
rect 880 25360 39200 25640
rect 800 13944 39200 25360
rect 800 13664 39120 13944
rect 800 2143 39200 13664
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< obsm4 >>
rect 19379 9011 19488 154597
rect 19968 9011 24781 154597
<< labels >>
rlabel metal3 s 39200 13744 40000 13864 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 275000 800 275120 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 125264 800 125384 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 88408 40000 88528 6 io_in[1]
port 4 nsew signal input
rlabel metal3 s 39200 163072 40000 163192 6 io_in[2]
port 5 nsew signal input
rlabel metal3 s 39200 237736 40000 237856 6 io_in[3]
port 6 nsew signal input
rlabel metal3 s 39200 312400 40000 312520 6 io_in[4]
port 7 nsew signal input
rlabel metal3 s 39200 387064 40000 387184 6 io_in[5]
port 8 nsew signal input
rlabel metal3 s 39200 461728 40000 461848 6 io_in[6]
port 9 nsew signal input
rlabel metal3 s 39200 536392 40000 536512 6 io_in[7]
port 10 nsew signal input
rlabel metal3 s 0 574472 800 574592 6 io_in[8]
port 11 nsew signal input
rlabel metal3 s 0 424736 800 424856 6 io_in[9]
port 12 nsew signal input
rlabel metal3 s 39200 63520 40000 63640 6 io_oeb[0]
port 13 nsew signal output
rlabel metal3 s 0 175176 800 175296 6 io_oeb[10]
port 14 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 io_oeb[11]
port 15 nsew signal output
rlabel metal3 s 39200 138184 40000 138304 6 io_oeb[1]
port 16 nsew signal output
rlabel metal3 s 39200 212848 40000 212968 6 io_oeb[2]
port 17 nsew signal output
rlabel metal3 s 39200 287512 40000 287632 6 io_oeb[3]
port 18 nsew signal output
rlabel metal3 s 39200 362176 40000 362296 6 io_oeb[4]
port 19 nsew signal output
rlabel metal3 s 39200 436840 40000 436960 6 io_oeb[5]
port 20 nsew signal output
rlabel metal3 s 39200 511504 40000 511624 6 io_oeb[6]
port 21 nsew signal output
rlabel metal3 s 39200 586168 40000 586288 6 io_oeb[7]
port 22 nsew signal output
rlabel metal3 s 0 474648 800 474768 6 io_oeb[8]
port 23 nsew signal output
rlabel metal3 s 0 324912 800 325032 6 io_oeb[9]
port 24 nsew signal output
rlabel metal3 s 39200 38632 40000 38752 6 io_out[0]
port 25 nsew signal output
rlabel metal3 s 0 225088 800 225208 6 io_out[10]
port 26 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 io_out[11]
port 27 nsew signal output
rlabel metal3 s 39200 113296 40000 113416 6 io_out[1]
port 28 nsew signal output
rlabel metal3 s 39200 187960 40000 188080 6 io_out[2]
port 29 nsew signal output
rlabel metal3 s 39200 262624 40000 262744 6 io_out[3]
port 30 nsew signal output
rlabel metal3 s 39200 337288 40000 337408 6 io_out[4]
port 31 nsew signal output
rlabel metal3 s 39200 411952 40000 412072 6 io_out[5]
port 32 nsew signal output
rlabel metal3 s 39200 486616 40000 486736 6 io_out[6]
port 33 nsew signal output
rlabel metal3 s 39200 561280 40000 561400 6 io_out[7]
port 34 nsew signal output
rlabel metal3 s 0 524560 800 524680 6 io_out[8]
port 35 nsew signal output
rlabel metal3 s 0 374824 800 374944 6 io_out[9]
port 36 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 38 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 39 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 40 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7734100
string GDS_FILE /home/hosni/OpenLane-tutorial/7-segment/openlane/user_proj_example1/runs/23_06_21_07_08/results/signoff/user_proj_example1.magic.gds
string GDS_START 565368
<< end >>


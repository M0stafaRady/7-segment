VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example1
  CLASS BLOCK ;
  FOREIGN user_proj_example1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.720 200.000 69.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.000 4.000 1375.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 626.320 4.000 626.920 ;
    END
  END io_in[11]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 442.040 200.000 442.640 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 815.360 200.000 815.960 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1188.680 200.000 1189.280 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1562.000 200.000 1562.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1935.320 200.000 1935.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2308.640 200.000 2309.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2681.960 200.000 2682.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2872.360 4.000 2872.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2123.680 4.000 2124.280 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 317.600 200.000 318.200 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 690.920 200.000 691.520 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1064.240 200.000 1064.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1437.560 200.000 1438.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1810.880 200.000 1811.480 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2184.200 200.000 2184.800 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2557.520 200.000 2558.120 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2930.840 200.000 2931.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2373.240 4.000 2373.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1624.560 4.000 1625.160 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.160 200.000 193.760 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_out[11]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 566.480 200.000 567.080 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 939.800 200.000 940.400 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1313.120 200.000 1313.720 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1686.440 200.000 1687.040 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2059.760 200.000 2060.360 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2433.080 200.000 2433.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2806.400 200.000 2807.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2622.800 4.000 2623.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1874.120 4.000 1874.720 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 195.430 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 195.410 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 195.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 2931.840 196.000 2986.725 ;
        RECT 4.000 2930.440 195.600 2931.840 ;
        RECT 4.000 2873.360 196.000 2930.440 ;
        RECT 4.400 2871.960 196.000 2873.360 ;
        RECT 4.000 2807.400 196.000 2871.960 ;
        RECT 4.000 2806.000 195.600 2807.400 ;
        RECT 4.000 2682.960 196.000 2806.000 ;
        RECT 4.000 2681.560 195.600 2682.960 ;
        RECT 4.000 2623.800 196.000 2681.560 ;
        RECT 4.400 2622.400 196.000 2623.800 ;
        RECT 4.000 2558.520 196.000 2622.400 ;
        RECT 4.000 2557.120 195.600 2558.520 ;
        RECT 4.000 2434.080 196.000 2557.120 ;
        RECT 4.000 2432.680 195.600 2434.080 ;
        RECT 4.000 2374.240 196.000 2432.680 ;
        RECT 4.400 2372.840 196.000 2374.240 ;
        RECT 4.000 2309.640 196.000 2372.840 ;
        RECT 4.000 2308.240 195.600 2309.640 ;
        RECT 4.000 2185.200 196.000 2308.240 ;
        RECT 4.000 2183.800 195.600 2185.200 ;
        RECT 4.000 2124.680 196.000 2183.800 ;
        RECT 4.400 2123.280 196.000 2124.680 ;
        RECT 4.000 2060.760 196.000 2123.280 ;
        RECT 4.000 2059.360 195.600 2060.760 ;
        RECT 4.000 1936.320 196.000 2059.360 ;
        RECT 4.000 1934.920 195.600 1936.320 ;
        RECT 4.000 1875.120 196.000 1934.920 ;
        RECT 4.400 1873.720 196.000 1875.120 ;
        RECT 4.000 1811.880 196.000 1873.720 ;
        RECT 4.000 1810.480 195.600 1811.880 ;
        RECT 4.000 1687.440 196.000 1810.480 ;
        RECT 4.000 1686.040 195.600 1687.440 ;
        RECT 4.000 1625.560 196.000 1686.040 ;
        RECT 4.400 1624.160 196.000 1625.560 ;
        RECT 4.000 1563.000 196.000 1624.160 ;
        RECT 4.000 1561.600 195.600 1563.000 ;
        RECT 4.000 1438.560 196.000 1561.600 ;
        RECT 4.000 1437.160 195.600 1438.560 ;
        RECT 4.000 1376.000 196.000 1437.160 ;
        RECT 4.400 1374.600 196.000 1376.000 ;
        RECT 4.000 1314.120 196.000 1374.600 ;
        RECT 4.000 1312.720 195.600 1314.120 ;
        RECT 4.000 1189.680 196.000 1312.720 ;
        RECT 4.000 1188.280 195.600 1189.680 ;
        RECT 4.000 1126.440 196.000 1188.280 ;
        RECT 4.400 1125.040 196.000 1126.440 ;
        RECT 4.000 1065.240 196.000 1125.040 ;
        RECT 4.000 1063.840 195.600 1065.240 ;
        RECT 4.000 940.800 196.000 1063.840 ;
        RECT 4.000 939.400 195.600 940.800 ;
        RECT 4.000 876.880 196.000 939.400 ;
        RECT 4.400 875.480 196.000 876.880 ;
        RECT 4.000 816.360 196.000 875.480 ;
        RECT 4.000 814.960 195.600 816.360 ;
        RECT 4.000 691.920 196.000 814.960 ;
        RECT 4.000 690.520 195.600 691.920 ;
        RECT 4.000 627.320 196.000 690.520 ;
        RECT 4.400 625.920 196.000 627.320 ;
        RECT 4.000 567.480 196.000 625.920 ;
        RECT 4.000 566.080 195.600 567.480 ;
        RECT 4.000 443.040 196.000 566.080 ;
        RECT 4.000 441.640 195.600 443.040 ;
        RECT 4.000 377.760 196.000 441.640 ;
        RECT 4.400 376.360 196.000 377.760 ;
        RECT 4.000 318.600 196.000 376.360 ;
        RECT 4.000 317.200 195.600 318.600 ;
        RECT 4.000 194.160 196.000 317.200 ;
        RECT 4.000 192.760 195.600 194.160 ;
        RECT 4.000 128.200 196.000 192.760 ;
        RECT 4.400 126.800 196.000 128.200 ;
        RECT 4.000 69.720 196.000 126.800 ;
        RECT 4.000 68.320 195.600 69.720 ;
        RECT 4.000 10.715 196.000 68.320 ;
      LAYER met4 ;
        RECT 96.895 45.055 97.440 772.985 ;
        RECT 99.840 45.055 123.905 772.985 ;
  END
END user_proj_example1
END LIBRARY

